library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROMWAV is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROMWAV is
	type rom is array(0 to  49151) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7C",X"7C",X"7B",X"7C",X"7B",X"C2",X"C2",X"84",X"7F",X"78",X"7B",X"78",X"7B",X"79",X"7B",X"7A",
		X"7A",X"7B",X"7A",X"7C",X"79",X"7B",X"76",X"AB",X"DF",X"E1",X"E5",X"E3",X"E4",X"E3",X"E4",X"E2",
		X"E2",X"E0",X"E0",X"DE",X"DF",X"DC",X"DF",X"D0",X"8B",X"74",X"71",X"6F",X"6F",X"6F",X"6F",X"6E",
		X"6F",X"6F",X"70",X"6F",X"70",X"6F",X"71",X"6F",X"AE",X"D7",X"D8",X"DB",X"D9",X"DA",X"D8",X"D9",
		X"D7",X"D8",X"D6",X"D8",X"D5",X"D7",X"D3",X"D7",X"9F",X"6D",X"6A",X"66",X"67",X"66",X"67",X"66",
		X"67",X"67",X"67",X"66",X"67",X"66",X"68",X"66",X"A4",X"CF",X"D0",X"D4",X"D1",X"D2",X"D1",X"D1",
		X"D0",X"CF",X"CF",X"CE",X"CF",X"CC",X"CF",X"C3",X"7F",X"63",X"62",X"5F",X"61",X"5E",X"60",X"5F",
		X"60",X"60",X"60",X"61",X"5F",X"62",X"5C",X"89",X"C4",X"C9",X"CE",X"CC",X"CD",X"CC",X"CB",X"CB",
		X"C9",X"CA",X"C7",X"C9",X"C5",X"CA",X"B6",X"72",X"5C",X"5B",X"59",X"5B",X"59",X"5B",X"59",X"5B",
		X"59",X"5B",X"59",X"5C",X"59",X"62",X"A4",X"C4",X"C4",X"C8",X"C5",X"C7",X"C4",X"C6",X"C4",X"C6",
		X"C3",X"C5",X"C3",X"C4",X"BE",X"7B",X"58",X"57",X"53",X"56",X"53",X"56",X"54",X"56",X"55",X"56",
		X"54",X"57",X"54",X"5F",X"A3",X"C0",X"C1",X"C4",X"C1",X"C2",X"C0",X"C2",X"BF",X"C1",X"BE",X"C1",
		X"BD",X"C3",X"A9",X"65",X"55",X"52",X"51",X"51",X"51",X"52",X"51",X"52",X"51",X"53",X"51",X"55",
		X"4F",X"85",X"B9",X"BB",X"C1",X"BE",X"C0",X"BE",X"BF",X"BD",X"BF",X"BC",X"BE",X"BB",X"BE",X"AC",
		X"66",X"51",X"4E",X"4D",X"4E",X"4D",X"4F",X"4E",X"4F",X"4E",X"50",X"4E",X"51",X"4F",X"8B",X"B8",
		X"B9",X"BE",X"BB",X"BD",X"BA",X"BC",X"B9",X"BB",X"B8",X"BB",X"B6",X"BE",X"93",X"56",X"50",X"4B",
		X"4D",X"4B",X"4D",X"4C",X"4E",X"4C",X"4E",X"4C",X"50",X"4A",X"69",X"AC",X"B6",X"BB",X"B9",X"BB",
		X"B9",X"BB",X"B9",X"BA",X"B8",X"BA",X"B6",X"BB",X"9F",X"5A",X"4D",X"49",X"4A",X"48",X"4A",X"49",
		X"4B",X"49",X"4C",X"49",X"4E",X"47",X"67",X"AB",X"B5",X"B9",X"B7",X"B9",X"B7",X"B8",X"B6",X"B8",
		X"B5",X"B8",X"B3",X"BA",X"8E",X"52",X"4C",X"48",X"49",X"48",X"49",X"49",X"4A",X"49",X"4B",X"4A",
		X"4C",X"4A",X"87",X"B3",X"B5",X"B8",X"B7",X"B7",X"B7",X"B6",X"B7",X"B5",X"B7",X"B4",X"B8",X"A9",
		X"63",X"4A",X"48",X"46",X"47",X"47",X"48",X"48",X"48",X"49",X"47",X"4B",X"45",X"74",X"AE",X"B2",
		X"B7",X"B6",X"B6",X"B6",X"B5",X"B5",X"B3",X"B4",X"B1",X"B5",X"A9",X"65",X"48",X"48",X"44",X"47",
		X"45",X"48",X"47",X"48",X"48",X"48",X"4A",X"46",X"7A",X"B0",X"B2",X"B7",X"B5",X"B6",X"B5",X"B4",
		X"B5",X"B3",X"B6",X"B1",X"B8",X"9B",X"58",X"4A",X"47",X"46",X"48",X"45",X"48",X"46",X"49",X"46",
		X"4A",X"45",X"54",X"98",X"B3",X"B3",X"B7",X"B4",X"B6",X"B3",X"B6",X"B3",X"B5",X"B3",X"B5",X"AE",
		X"6D",X"48",X"48",X"43",X"47",X"44",X"47",X"45",X"47",X"46",X"48",X"48",X"49",X"88",X"B2",X"B2",
		X"B7",X"B4",X"B6",X"B3",X"B4",X"B3",X"B3",X"B3",X"B2",X"B2",X"76",X"49",X"49",X"44",X"47",X"45",
		X"47",X"46",X"47",X"47",X"48",X"48",X"49",X"87",X"B1",X"B1",X"B6",X"B3",X"B5",X"B2",X"B4",X"B2",
		X"B3",X"B2",X"B3",X"AF",X"6E",X"49",X"49",X"44",X"47",X"44",X"47",X"45",X"47",X"45",X"48",X"44",
		X"52",X"98",X"B2",X"B2",X"B5",X"B3",X"B5",X"B3",X"B5",X"B2",X"B6",X"B1",X"B8",X"9B",X"57",X"49",
		X"45",X"45",X"46",X"45",X"47",X"46",X"48",X"46",X"4A",X"44",X"77",X"AF",X"B2",X"B7",X"B4",X"B6",
		X"B5",X"B6",X"B4",X"B4",X"B2",X"B3",X"AE",X"6B",X"49",X"48",X"44",X"47",X"45",X"48",X"45",X"48",
		X"45",X"4A",X"43",X"62",X"A6",X"B1",X"B5",X"B4",X"B4",X"B4",X"B4",X"B3",X"B2",X"B2",X"B0",X"B2",
		X"76",X"48",X"48",X"43",X"46",X"44",X"47",X"45",X"48",X"45",X"4A",X"44",X"5D",X"A3",X"B1",X"B5",
		X"B5",X"B4",X"B4",X"B4",X"B4",X"B3",X"B4",X"B3",X"B4",X"77",X"4B",X"4A",X"45",X"48",X"46",X"49",
		X"46",X"49",X"46",X"4A",X"45",X"5C",X"A2",X"B2",X"B5",X"B6",X"B5",X"B7",X"B5",X"B7",X"B4",X"B7",
		X"B2",X"BA",X"96",X"55",X"49",X"46",X"45",X"47",X"45",X"48",X"45",X"49",X"45",X"4B",X"44",X"62",
		X"A5",X"B4",X"B6",X"B7",X"B6",X"B7",X"B5",X"B6",X"B3",X"B3",X"B3",X"B3",X"AF",X"6F",X"4A",X"48",
		X"46",X"47",X"47",X"48",X"48",X"48",X"49",X"48",X"4B",X"47",X"5A",X"A0",X"B2",X"B6",X"B5",X"B6",
		X"B4",X"B6",X"B3",X"B7",X"9D",X"5A",X"4D",X"49",X"49",X"48",X"4A",X"49",X"4A",X"4A",X"4A",X"4B",
		X"4A",X"4B",X"4B",X"4C",X"4C",X"4D",X"4D",X"4E",X"4E",X"4F",X"4F",X"50",X"4F",X"50",X"50",X"50",
		X"50",X"50",X"50",X"50",X"51",X"51",X"52",X"52",X"52",X"52",X"53",X"53",X"54",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"56",X"56",X"56",X"56",X"57",X"57",X"57",X"58",X"58",X"59",X"59",X"59",
		X"5A",X"5A",X"5A",X"5A",X"5A",X"5B",X"5B",X"5B",X"5B",X"5B",X"5B",X"5C",X"5C",X"5C",X"5D",X"5D",
		X"5D",X"5D",X"5D",X"5D",X"5D",X"5E",X"5E",X"5E",X"5E",X"5F",X"5F",X"5F",X"5F",X"60",X"60",X"60",
		X"61",X"61",X"61",X"61",X"62",X"62",X"62",X"62",X"63",X"63",X"63",X"63",X"63",X"64",X"64",X"64",
		X"64",X"64",X"65",X"65",X"65",X"65",X"66",X"66",X"66",X"66",X"66",X"67",X"67",X"67",X"67",X"67",
		X"67",X"67",X"68",X"68",X"68",X"68",X"68",X"68",X"69",X"69",X"69",X"69",X"69",X"69",X"6A",X"6A",
		X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",
		X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6F",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",
		X"71",X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"73",X"73",X"73",
		X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"75",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",
		X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"78",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",X"78",
		X"78",X"78",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"80",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7B",X"7C",X"7A",X"7D",X"77",X"9A",X"D6",X"A4",X"81",X"7D",X"79",X"7B",X"79",X"7B",X"79",X"7B",
		X"79",X"7C",X"79",X"7C",X"79",X"7C",X"78",X"7C",X"75",X"96",X"D3",X"DE",X"E3",X"E2",X"E3",X"E1",
		X"E2",X"E1",X"E1",X"E0",X"E0",X"DD",X"DF",X"DC",X"DE",X"DA",X"DE",X"CB",X"89",X"75",X"71",X"70",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"70",X"6F",X"71",X"6E",X"72",X"6D",X"84",X"C5",X"D6",
		X"D8",X"D9",X"D8",X"D8",X"D7",X"D7",X"D6",X"D6",X"D6",X"D6",X"D6",X"D4",X"D6",X"D2",X"D6",X"AD",
		X"73",X"6B",X"66",X"67",X"66",X"67",X"67",X"67",X"67",X"67",X"68",X"66",X"68",X"66",X"69",X"65",
		X"70",X"B0",X"CE",X"CF",X"D2",X"D0",X"D2",X"CF",X"D0",X"CE",X"CF",X"CD",X"CE",X"CD",X"CD",X"CD",
		X"CB",X"CD",X"97",X"68",X"65",X"5F",X"61",X"5F",X"60",X"5F",X"60",X"60",X"60",X"60",X"60",X"61",
		X"60",X"62",X"5E",X"91",X"C3",X"C7",X"CC",X"CA",X"CC",X"CA",X"CB",X"CA",X"C9",X"C8",X"C8",X"C7",
		X"C6",X"C7",X"C5",X"C6",X"8F",X"61",X"5E",X"59",X"5B",X"59",X"5B",X"5A",X"5B",X"5A",X"5B",X"5A",
		X"5C",X"5A",X"5C",X"59",X"64",X"A6",X"C1",X"C4",X"C6",X"C4",X"C5",X"C4",X"C5",X"C3",X"C5",X"C3",
		X"C4",X"C2",X"C4",X"C0",X"C6",X"9D",X"62",X"5A",X"54",X"56",X"54",X"56",X"55",X"56",X"55",X"57",
		X"56",X"57",X"56",X"57",X"55",X"62",X"A5",X"BD",X"C0",X"C2",X"C1",X"C1",X"C0",X"C0",X"BF",X"BF",
		X"BF",X"BF",X"BE",X"BF",X"BD",X"BC",X"7F",X"59",X"55",X"51",X"53",X"51",X"53",X"52",X"53",X"52",
		X"53",X"52",X"54",X"52",X"55",X"53",X"8D",X"B7",X"BB",X"BF",X"BD",X"BE",X"BD",X"BE",X"BD",X"BD",
		X"BC",X"BD",X"BB",X"BC",X"B9",X"B9",X"7D",X"55",X"51",X"4E",X"4F",X"4E",X"4F",X"4F",X"4F",X"50",
		X"4F",X"50",X"50",X"51",X"4F",X"58",X"99",X"B7",X"BA",X"BC",X"BA",X"BB",X"BA",X"BA",X"BA",X"B9",
		X"BA",X"B8",X"BA",X"B6",X"BC",X"A1",X"60",X"51",X"4D",X"4D",X"4D",X"4D",X"4E",X"4D",X"4E",X"4D",
		X"4E",X"4E",X"4E",X"4F",X"4E",X"84",X"B3",X"B5",X"BA",X"B8",X"BA",X"B9",X"B9",X"B9",X"B8",X"B9",
		X"B7",X"B9",X"B5",X"BA",X"9F",X"5F",X"4E",X"4B",X"4A",X"4B",X"4A",X"4C",X"4A",X"4C",X"4A",X"4D",
		X"4B",X"4D",X"4B",X"52",X"91",X"B3",X"B4",X"B9",X"B6",X"B8",X"B5",X"B7",X"B5",X"B6",X"B5",X"B5",
		X"B5",X"B3",X"B5",X"81",X"51",X"4D",X"48",X"4B",X"49",X"4A",X"4A",X"4B",X"4B",X"4B",X"4C",X"4A",
		X"4E",X"49",X"78",X"AE",X"B2",X"B7",X"B6",X"B7",X"B6",X"B6",X"B6",X"B5",X"B6",X"B4",X"B6",X"B2",
		X"B8",X"8A",X"53",X"4C",X"47",X"49",X"47",X"48",X"48",X"49",X"49",X"49",X"4A",X"49",X"4B",X"48",
		X"7B",X"AD",X"B1",X"B6",X"B4",X"B6",X"B4",X"B5",X"B3",X"B3",X"B2",X"B2",X"B2",X"B1",X"B1",X"77",
		X"4D",X"4A",X"45",X"48",X"46",X"49",X"47",X"49",X"48",X"4A",X"48",X"4B",X"48",X"54",X"96",X"B0",
		X"B3",X"B6",X"B4",X"B5",X"B3",X"B5",X"B3",X"B5",X"B2",X"B5",X"B1",X"B7",X"95",X"57",X"4C",X"47",
		X"48",X"47",X"48",X"48",X"48",X"48",X"48",X"49",X"49",X"4A",X"4B",X"87",X"AF",X"B1",X"B5",X"B3",
		X"B5",X"B3",X"B5",X"B3",X"B5",X"B2",X"B5",X"B0",X"B7",X"96",X"56",X"4B",X"46",X"47",X"46",X"47",
		X"46",X"48",X"47",X"48",X"48",X"49",X"48",X"4F",X"90",X"AF",X"B2",X"B5",X"B4",X"B5",X"B3",X"B4",
		X"B2",X"B3",X"B1",X"B3",X"AF",X"B4",X"83",X"4F",X"4A",X"45",X"48",X"46",X"48",X"46",X"49",X"47",
		X"49",X"47",X"4B",X"44",X"64",X"A4",X"AF",X"B4",X"B3",X"B4",X"B2",X"B3",X"B2",X"B3",X"B1",X"B3",
		X"B0",X"B4",X"A3",X"60",X"4C",X"47",X"47",X"46",X"47",X"47",X"47",X"47",X"47",X"47",X"48",X"46",
		X"51",X"95",X"AE",X"B2",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"B3",X"AC",X"6A",
		X"4C",X"48",X"46",X"47",X"46",X"47",X"47",X"47",X"48",X"48",X"49",X"48",X"50",X"94",X"AF",X"B3",
		X"B5",X"B5",X"B4",X"B5",X"B4",X"B4",X"B3",X"B3",X"B1",X"B3",X"A7",X"63",X"4C",X"47",X"47",X"46",
		X"47",X"47",X"48",X"47",X"49",X"47",X"4A",X"45",X"5B",X"9E",X"AF",X"B4",X"B3",X"B4",X"B3",X"B4",
		X"B2",X"B3",X"B0",X"B2",X"AE",X"B4",X"92",X"54",X"4A",X"45",X"46",X"45",X"47",X"46",X"48",X"47",
		X"49",X"47",X"4A",X"46",X"79",X"AB",X"B0",X"B5",X"B3",X"B4",X"B3",X"B3",X"B2",X"B3",X"B2",X"B3",
		X"B3",X"AE",X"6F",X"4E",X"4B",X"47",X"49",X"48",X"49",X"48",X"49",X"49",X"49",X"4A",X"48",X"56",
		X"99",X"AF",X"B4",X"B4",X"B5",X"B5",X"B5",X"B5",X"B4",X"B5",X"B4",X"B4",X"B5",X"AE",X"6C",X"4D",
		X"49",X"46",X"47",X"46",X"48",X"47",X"48",X"47",X"4A",X"47",X"4C",X"46",X"75",X"AC",X"B1",X"B6",
		X"B4",X"B6",X"B5",X"B6",X"B4",X"B4",X"B2",X"B2",X"B2",X"B1",X"AF",X"76",X"4D",X"4A",X"46",X"49",
		X"47",X"49",X"48",X"4A",X"49",X"49",X"49",X"4B",X"4B",X"4B",X"82",X"AE",X"B1",X"B6",X"B3",X"B5",
		X"B3",X"B4",X"B3",X"B3",X"B0",X"74",X"50",X"4D",X"49",X"4B",X"49",X"4B",X"4A",X"4B",X"4A",X"4B",
		X"4B",X"4B",X"4B",X"4C",X"4D",X"4D",X"4D",X"4E",X"4E",X"4F",X"4F",X"50",X"50",X"50",X"50",X"50",
		X"51",X"50",X"51",X"51",X"51",X"51",X"51",X"51",X"52",X"52",X"52",X"52",X"53",X"53",X"54",X"54",
		X"54",X"55",X"55",X"56",X"56",X"56",X"56",X"56",X"56",X"56",X"57",X"57",X"57",X"57",X"58",X"58",
		X"58",X"59",X"59",X"59",X"5A",X"5A",X"5A",X"5B",X"5B",X"5B",X"5B",X"5B",X"5B",X"5B",X"5C",X"5C",
		X"5C",X"5C",X"5C",X"5D",X"5D",X"5D",X"5D",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5F",X"5F",
		X"5F",X"5F",X"5F",X"5F",X"60",X"60",X"60",X"61",X"61",X"61",X"61",X"62",X"62",X"62",X"62",X"63",
		X"63",X"63",X"63",X"63",X"64",X"64",X"64",X"64",X"64",X"64",X"64",X"65",X"65",X"65",X"65",X"65",
		X"66",X"66",X"66",X"66",X"66",X"66",X"67",X"67",X"67",X"67",X"67",X"68",X"68",X"68",X"68",X"68",
		X"68",X"68",X"68",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"6A",X"6A",X"6A",X"6A",X"6A",X"6B",
		X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",
		X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6F",X"6F",X"6F",X"6F",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"73",X"73",X"73",
		X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",
		X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"80",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7D",X"7B",X"7C",X"7B",X"7C",X"7B",X"B4",X"D4",X"9C",X"83",X"7C",X"7A",X"7A",X"79",X"7A",X"79",
		X"7A",X"7A",X"7B",X"7A",X"7B",X"7A",X"7B",X"7A",X"7C",X"79",X"7B",X"76",X"8A",X"C9",X"DC",X"E1",
		X"E2",X"E2",X"E2",X"E2",X"E2",X"E1",X"E1",X"E0",X"E0",X"DE",X"DE",X"DD",X"DE",X"DC",X"DD",X"DA",
		X"DD",X"AB",X"7C",X"75",X"70",X"71",X"6F",X"70",X"6F",X"70",X"6F",X"70",X"6F",X"70",X"6F",X"70",
		X"6F",X"71",X"6E",X"72",X"6C",X"91",X"CA",X"D4",X"D9",X"D8",X"D9",X"D8",X"D8",X"D7",X"D7",X"D6",
		X"D6",X"D6",X"D6",X"D5",X"D6",X"D4",X"D6",X"D2",X"D6",X"B0",X"78",X"6D",X"67",X"67",X"66",X"67",
		X"67",X"67",X"67",X"67",X"67",X"67",X"67",X"67",X"67",X"67",X"67",X"68",X"68",X"9D",X"C9",X"CD",
		X"D2",X"D0",X"D2",X"D0",X"D1",X"CF",X"CF",X"CF",X"CE",X"CE",X"CD",X"CE",X"CC",X"CE",X"CA",X"CF",
		X"B7",X"7A",X"67",X"62",X"60",X"61",X"60",X"60",X"5F",X"61",X"5F",X"61",X"5F",X"61",X"60",X"62",
		X"60",X"62",X"5F",X"69",X"A6",X"C5",X"C8",X"CC",X"CA",X"CC",X"CA",X"CB",X"CA",X"CB",X"C8",X"C9",
		X"C7",X"C8",X"C6",X"C7",X"C5",X"C7",X"C0",X"84",X"62",X"5E",X"5A",X"5B",X"5A",X"5B",X"5A",X"5B",
		X"5A",X"5B",X"5A",X"5C",X"5A",X"5C",X"5A",X"5C",X"59",X"68",X"A7",X"BF",X"C4",X"C6",X"C5",X"C5",
		X"C4",X"C5",X"C4",X"C5",X"C3",X"C4",X"C3",X"C4",X"C2",X"C4",X"C0",X"C5",X"9F",X"66",X"5B",X"55",
		X"56",X"54",X"56",X"55",X"56",X"55",X"56",X"56",X"57",X"56",X"56",X"56",X"57",X"56",X"5D",X"9B",
		X"BA",X"BF",X"C2",X"C1",X"C1",X"C0",X"C1",X"BF",X"C0",X"BF",X"C0",X"BE",X"BF",X"BD",X"BF",X"BC",
		X"C0",X"8E",X"5F",X"57",X"52",X"53",X"51",X"53",X"52",X"53",X"52",X"53",X"52",X"53",X"52",X"54",
		X"52",X"56",X"50",X"7B",X"B0",X"B9",X"BE",X"BD",X"BF",X"BD",X"BE",X"BD",X"BE",X"BD",X"BD",X"BC",
		X"BD",X"BB",X"BD",X"B8",X"BD",X"91",X"5C",X"53",X"4E",X"4F",X"4E",X"4F",X"4E",X"4F",X"4F",X"4F",
		X"50",X"50",X"50",X"50",X"50",X"51",X"50",X"84",X"B2",X"B7",X"BC",X"BA",X"BC",X"BA",X"BB",X"BA",
		X"BA",X"BA",X"B9",X"B9",X"B8",X"B9",X"B7",X"BA",X"AF",X"73",X"56",X"52",X"4F",X"51",X"4F",X"51",
		X"51",X"52",X"4F",X"4E",X"4E",X"4D",X"4E",X"4D",X"50",X"4B",X"6F",X"A4",X"AC",X"B1",X"B0",X"B1",
		X"B0",X"B1",X"B7",X"B7",X"B8",X"B7",X"B8",X"B6",X"B8",X"B5",X"B8",X"AB",X"75",X"5C",X"59",X"56",
		X"58",X"52",X"4D",X"4A",X"4B",X"4A",X"4B",X"4A",X"4B",X"4B",X"4C",X"4C",X"4C",X"7A",X"9E",X"A1",
		X"A6",X"AE",X"B6",X"B5",X"B7",X"B5",X"B6",X"B5",X"B5",X"B5",X"B4",X"B5",X"B2",X"B6",X"91",X"6A",
		X"5E",X"4D",X"4A",X"48",X"49",X"49",X"49",X"4A",X"49",X"4A",X"4A",X"4B",X"4A",X"4C",X"49",X"6A",
		X"9F",X"B0",X"B5",X"B5",X"B6",X"B5",X"B5",X"B5",X"B5",X"B5",X"B5",X"B4",X"B4",X"B4",X"B4",X"AE",
		X"7B",X"53",X"4C",X"47",X"49",X"47",X"49",X"48",X"49",X"48",X"49",X"49",X"49",X"4A",X"49",X"5C",
		X"6C",X"94",X"B0",X"B2",X"B6",X"B4",X"B6",X"B4",X"B5",X"B4",X"B5",X"B3",X"B4",X"B2",X"B3",X"9B",
		X"8D",X"83",X"5B",X"4B",X"48",X"47",X"47",X"47",X"47",X"48",X"48",X"48",X"49",X"49",X"49",X"5B",
		X"74",X"74",X"8C",X"AB",X"B2",X"B5",X"B5",X"B5",X"B5",X"B4",X"B4",X"B3",X"B3",X"B3",X"B3",X"AF",
		X"93",X"83",X"7E",X"5D",X"4C",X"49",X"48",X"48",X"48",X"48",X"48",X"49",X"48",X"49",X"49",X"4A",
		X"4D",X"6E",X"7C",X"92",X"AE",X"B1",X"B5",X"B3",X"B5",X"B3",X"B5",X"B2",X"B4",X"98",X"7F",X"7B",
		X"79",X"78",X"78",X"70",X"54",X"4C",X"49",X"49",X"48",X"49",X"49",X"4A",X"49",X"4A",X"4B",X"4B",
		X"4B",X"4C",X"4C",X"4E",X"67",X"73",X"75",X"76",X"76",X"76",X"75",X"75",X"74",X"74",X"74",X"74",
		X"73",X"73",X"72",X"72",X"5F",X"51",X"4F",X"4E",X"4F",X"4F",X"4F",X"4F",X"50",X"50",X"51",X"51",
		X"52",X"51",X"52",X"52",X"62",X"6F",X"70",X"72",X"71",X"71",X"71",X"71",X"70",X"71",X"70",X"70",
		X"70",X"70",X"70",X"70",X"63",X"58",X"56",X"55",X"56",X"56",X"56",X"56",X"56",X"56",X"57",X"57",
		X"57",X"57",X"58",X"58",X"64",X"6D",X"6E",X"6F",X"6E",X"6F",X"6F",X"6E",X"6E",X"6E",X"6D",X"6D",
		X"6D",X"6D",X"6E",X"6C",X"62",X"5C",X"5C",X"5B",X"5C",X"5C",X"5D",X"5D",X"5D",X"5E",X"5E",X"5E",
		X"5E",X"5F",X"5F",X"62",X"6A",X"6C",X"6C",X"6D",X"6D",X"6D",X"6D",X"6C",X"6C",X"6C",X"6C",X"6C",
		X"6C",X"6C",X"6C",X"69",X"65",X"64",X"64",X"64",X"65",X"65",X"65",X"65",X"66",X"66",X"66",X"66",
		X"67",X"67",X"67",X"6A",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",
		X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",
		X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6F",X"6F",X"6F",X"6F",
		X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"71",X"71",
		X"71",X"71",X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"73",
		X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"74",
		X"74",X"74",X"74",X"75",X"74",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"76",
		X"76",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"79",
		X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",
		X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7C",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"81",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"80",X"81",X"81",X"80",X"80",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"9B",X"B9",X"B7",X"BF",X"B7",X"BF",X"CA",X"C7",X"CE",X"C8",X"BC",X"BF",X"B6",X"A9",X"B9",X"B6",
		X"BE",X"C6",X"BF",X"CA",X"CA",X"C0",X"C0",X"B8",X"B1",X"B9",X"A4",X"B0",X"A8",X"AF",X"B4",X"B3",
		X"B3",X"BA",X"B7",X"C0",X"B9",X"BB",X"C8",X"B6",X"CE",X"AD",X"C5",X"B3",X"BC",X"B8",X"AF",X"BB",
		X"AB",X"BC",X"A7",X"B6",X"AB",X"B2",X"B0",X"A8",X"B3",X"A7",X"B2",X"AC",X"A7",X"B5",X"A5",X"B8",
		X"AD",X"A9",X"BF",X"A3",X"C4",X"B0",X"A9",X"BF",X"A3",X"B3",X"A8",X"9E",X"A8",X"A3",X"93",X"A7",
		X"8B",X"91",X"A4",X"88",X"9D",X"A0",X"99",X"A5",X"B0",X"96",X"B6",X"B0",X"9B",X"A5",X"A1",X"8A",
		X"98",X"9C",X"81",X"96",X"A0",X"95",X"A0",X"B7",X"9C",X"99",X"A8",X"98",X"83",X"94",X"96",X"87",
		X"99",X"AC",X"9C",X"93",X"A6",X"9D",X"83",X"88",X"9B",X"91",X"8E",X"A8",X"B1",X"90",X"8A",X"97",
		X"94",X"80",X"89",X"A5",X"A5",X"8F",X"8F",X"98",X"8D",X"7E",X"8B",X"A9",X"A5",X"89",X"85",X"92",
		X"93",X"85",X"84",X"9C",X"A7",X"91",X"75",X"7D",X"96",X"9C",X"91",X"88",X"8D",X"91",X"8A",X"82",
		X"89",X"9A",X"9A",X"85",X"71",X"7F",X"9D",X"AC",X"91",X"75",X"72",X"91",X"A2",X"9C",X"81",X"75",
		X"81",X"97",X"9D",X"8B",X"7B",X"79",X"8C",X"97",X"99",X"81",X"7B",X"78",X"95",X"99",X"9A",X"7A",
		X"72",X"75",X"97",X"A2",X"98",X"77",X"65",X"78",X"90",X"A1",X"8D",X"85",X"6F",X"86",X"7D",X"96",
		X"7F",X"98",X"7D",X"8E",X"69",X"7D",X"7B",X"A2",X"A3",X"84",X"80",X"5F",X"8F",X"6D",X"A5",X"72",
		X"AE",X"73",X"94",X"57",X"6F",X"86",X"87",X"AC",X"6C",X"A7",X"60",X"A0",X"54",X"7E",X"7A",X"8B",
		X"B0",X"70",X"A8",X"67",X"91",X"64",X"5A",X"91",X"6C",X"AE",X"70",X"95",X"96",X"73",X"96",X"41",
		X"88",X"70",X"71",X"98",X"6A",X"C0",X"89",X"7C",X"97",X"5E",X"9B",X"53",X"59",X"90",X"5C",X"9F",
		X"78",X"89",X"C5",X"6C",X"95",X"85",X"68",X"9A",X"44",X"67",X"8D",X"52",X"92",X"7B",X"7A",X"B5",
		X"6D",X"8E",X"AE",X"6B",X"96",X"7E",X"5D",X"9A",X"4D",X"54",X"99",X"59",X"77",X"8F",X"62",X"9E",
		X"94",X"66",X"C3",X"98",X"68",X"A8",X"7C",X"71",X"9A",X"5D",X"66",X"97",X"40",X"5B",X"99",X"52",
		X"63",X"93",X"5D",X"75",X"9B",X"66",X"87",X"AB",X"65",X"89",X"C7",X"71",X"7C",X"BB",X"79",X"6D",
		X"A4",X"78",X"67",X"9B",X"71",X"59",X"93",X"71",X"47",X"8E",X"80",X"31",X"72",X"92",X"3C",X"58",
		X"9C",X"60",X"4F",X"92",X"79",X"4F",X"88",X"91",X"5C",X"7A",X"9C",X"69",X"6C",X"A4",X"82",X"62",
		X"9A",X"9C",X"5F",X"80",X"B3",X"7A",X"67",X"AD",X"A0",X"5C",X"8A",X"C0",X"7C",X"66",X"B5",X"AA",
		X"5B",X"84",X"C9",X"86",X"5D",X"AE",X"BB",X"63",X"72",X"C9",X"A0",X"59",X"97",X"C9",X"7C",X"5C",
		X"B1",X"BA",X"65",X"71",X"BD",X"9F",X"56",X"83",X"C0",X"8A",X"59",X"95",X"B5",X"75",X"5B",X"9F",
		X"AC",X"6A",X"64",X"9F",X"9B",X"5F",X"63",X"9B",X"95",X"5E",X"63",X"92",X"8E",X"57",X"5C",X"8F",
		X"90",X"54",X"54",X"86",X"8E",X"47",X"45",X"86",X"92",X"41",X"35",X"82",X"90",X"40",X"30",X"85",
		X"92",X"57",X"38",X"80",X"91",X"71",X"48",X"7A",X"9A",X"8C",X"53",X"6C",X"9D",X"A6",X"69",X"60",
		X"A5",X"C4",X"7E",X"52",X"98",X"C4",X"98",X"51",X"83",X"99",X"A7",X"51",X"67",X"74",X"AD",X"69",
		X"4F",X"50",X"97",X"8C",X"36",X"30",X"78",X"A9",X"54",X"4F",X"4B",X"B1",X"72",X"80",X"3D",X"9C",
		X"9D",X"A3",X"55",X"63",X"BD",X"BF",X"90",X"40",X"A5",X"8F",X"BE",X"40",X"77",X"63",X"B1",X"80",
		X"46",X"49",X"68",X"BA",X"48",X"57",X"31",X"B2",X"85",X"83",X"52",X"5F",X"B5",X"9A",X"A6",X"37",
		X"99",X"AE",X"C7",X"6C",X"4E",X"8E",X"84",X"BE",X"49",X"62",X"49",X"99",X"A0",X"40",X"47",X"40",
		X"BF",X"7A",X"84",X"4C",X"5F",X"B6",X"A6",X"B1",X"38",X"87",X"88",X"AD",X"96",X"3D",X"55",X"48",
		X"C2",X"7A",X"79",X"51",X"55",X"BE",X"B6",X"C2",X"41",X"74",X"58",X"97",X"A7",X"5A",X"6C",X"41",
		X"81",X"45",X"36",X"34",X"33",X"36",X"32",X"37",X"33",X"37",X"34",X"38",X"35",X"39",X"36",X"3A",
		X"38",X"3B",X"39",X"3C",X"3A",X"3C",X"3B",X"3C",X"3C",X"3D",X"3D",X"3D",X"3E",X"3E",X"3F",X"3F",
		X"40",X"40",X"41",X"41",X"42",X"42",X"43",X"43",X"43",X"43",X"44",X"44",X"45",X"45",X"46",X"46",
		X"47",X"47",X"48",X"49",X"49",X"4A",X"4A",X"4B",X"4B",X"4B",X"4B",X"4C",X"4C",X"4D",X"4D",X"4D",
		X"4E",X"4E",X"4E",X"4F",X"4F",X"50",X"50",X"50",X"51",X"51",X"51",X"51",X"51",X"51",X"52",X"52",
		X"52",X"53",X"53",X"54",X"54",X"54",X"55",X"56",X"56",X"57",X"57",X"57",X"57",X"58",X"58",X"58",
		X"59",X"59",X"59",X"5A",X"5A",X"5A",X"5A",X"5B",X"5B",X"5B",X"5C",X"5C",X"5C",X"5D",X"5D",X"5D",
		X"5D",X"5E",X"5E",X"5E",X"5E",X"5E",X"5F",X"5F",X"5F",X"5F",X"60",X"60",X"60",X"61",X"61",X"61",
		X"61",X"62",X"62",X"62",X"62",X"63",X"63",X"63",X"63",X"64",X"64",X"64",X"65",X"65",X"65",X"65",
		X"66",X"66",X"66",X"66",X"67",X"67",X"67",X"67",X"68",X"68",X"68",X"68",X"69",X"69",X"69",X"69",
		X"69",X"69",X"6A",X"6A",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",
		X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6E",
		X"6E",X"6E",X"6F",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"71",
		X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"73",X"73",X"73",X"73",X"73",X"73",
		X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",
		X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"76",
		X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"79",X"79",X"79",X"79",X"79",
		X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"82",X"82",X"82",
		X"82",X"81",X"82",X"81",X"82",X"81",X"82",X"82",X"82",X"82",X"81",X"82",X"82",X"81",X"81",X"82",
		X"82",X"81",X"81",X"82",X"82",X"82",X"82",X"81",X"82",X"82",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"82",X"81",X"81",X"81",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"81",X"81",X"80",X"80",
		X"9D",X"BA",X"B7",X"C0",X"BA",X"BA",X"C7",X"CA",X"C9",X"D0",X"C7",X"BD",X"BF",X"BC",X"A8",X"B8",
		X"B6",X"BC",X"C0",X"CA",X"BC",X"D0",X"C8",X"C2",X"C2",X"B9",X"B6",X"B3",X"B7",X"9E",X"BA",X"A0",
		X"B7",X"B2",X"B4",X"B5",X"B5",X"BF",X"B4",X"C9",X"AE",X"CA",X"BF",X"BB",X"CF",X"AE",X"C3",X"BA",
		X"B5",X"C3",X"AB",X"BC",X"B3",X"B2",X"BA",X"A9",X"B5",X"AF",X"AE",X"B6",X"A7",X"B0",X"B0",X"A7",
		X"B6",X"A9",X"A9",X"B6",X"A7",X"B3",X"B7",X"A1",X"BC",X"B3",X"A9",X"CA",X"A9",X"AD",X"C0",X"A5",
		X"AF",X"B0",X"9E",X"A4",X"AB",X"9B",X"98",X"A7",X"89",X"90",X"A7",X"8A",X"96",X"A3",X"9B",X"9C",
		X"AE",X"AA",X"98",X"BA",X"B1",X"9A",X"A6",X"A3",X"93",X"8A",X"A4",X"8F",X"83",X"9C",X"9E",X"98",
		X"9C",X"BA",X"A3",X"96",X"A5",X"A4",X"8F",X"82",X"9B",X"91",X"8A",X"95",X"AD",X"A3",X"90",X"A1",
		X"A4",X"96",X"7C",X"90",X"99",X"92",X"8E",X"A2",X"B8",X"97",X"8C",X"8C",X"9D",X"8B",X"80",X"8C",
		X"A6",X"A8",X"8F",X"91",X"92",X"9A",X"7F",X"84",X"91",X"B1",X"9F",X"8A",X"84",X"91",X"96",X"88",
		X"83",X"8C",X"A9",X"A0",X"8D",X"70",X"82",X"92",X"A1",X"91",X"8C",X"87",X"93",X"8D",X"88",X"80",
		X"8E",X"9A",X"9C",X"87",X"72",X"78",X"90",X"AC",X"A2",X"88",X"6D",X"7A",X"8E",X"A8",X"99",X"8C",
		X"6F",X"81",X"87",X"A5",X"90",X"8F",X"70",X"83",X"84",X"9E",X"95",X"8A",X"7D",X"71",X"8F",X"8A",
		X"AF",X"7E",X"93",X"55",X"90",X"77",X"B9",X"8F",X"8E",X"6B",X"5E",X"92",X"7D",X"BD",X"6F",X"A2",
		X"58",X"93",X"75",X"8E",X"93",X"79",X"A5",X"6A",X"9F",X"5B",X"82",X"7C",X"8C",X"BD",X"77",X"9D",
		X"58",X"7C",X"82",X"74",X"A8",X"6C",X"B0",X"7D",X"86",X"7F",X"45",X"93",X"6F",X"A4",X"9A",X"73",
		X"A4",X"67",X"92",X"75",X"56",X"95",X"69",X"AB",X"9D",X"75",X"A9",X"67",X"88",X"7B",X"43",X"91",
		X"72",X"8A",X"A6",X"66",X"A3",X"8E",X"73",X"9A",X"4B",X"6B",X"8F",X"57",X"96",X"81",X"79",X"C7",
		X"80",X"7C",X"9D",X"5E",X"8D",X"7B",X"38",X"85",X"79",X"65",X"A5",X"71",X"89",X"CA",X"77",X"81",
		X"9E",X"61",X"89",X"84",X"36",X"7B",X"86",X"52",X"8D",X"87",X"6B",X"AE",X"93",X"65",X"AF",X"98",
		X"6B",X"9B",X"7D",X"59",X"97",X"68",X"38",X"8D",X"7E",X"53",X"8C",X"84",X"63",X"A1",X"9A",X"61",
		X"AF",X"BB",X"65",X"8B",X"A4",X"6A",X"7D",X"99",X"5A",X"62",X"99",X"54",X"3D",X"92",X"79",X"45",
		X"7C",X"8C",X"57",X"79",X"9C",X"6A",X"77",X"AE",X"83",X"60",X"B6",X"B3",X"63",X"89",X"BB",X"7C",
		X"65",X"9F",X"8C",X"5F",X"85",X"97",X"5B",X"66",X"97",X"6B",X"46",X"85",X"91",X"3B",X"4C",X"98",
		X"6E",X"30",X"72",X"99",X"5A",X"4E",X"8D",X"86",X"4F",X"6E",X"9C",X"76",X"5B",X"8B",X"97",X"65",
		X"6B",X"A2",X"8D",X"61",X"82",X"AB",X"7C",X"5E",X"96",X"B0",X"72",X"67",X"A8",X"AD",X"66",X"6D",
		X"B7",X"AA",X"63",X"79",X"C1",X"A1",X"5B",X"7B",X"CA",X"9D",X"5D",X"83",X"CC",X"97",X"59",X"83",
		X"D1",X"9A",X"5C",X"86",X"CD",X"9B",X"57",X"81",X"C8",X"A3",X"57",X"7F",X"BB",X"AA",X"53",X"77",
		X"B0",X"B5",X"5A",X"72",X"A1",X"B7",X"62",X"64",X"97",X"B6",X"76",X"5A",X"8C",X"A3",X"8B",X"48",
		X"7F",X"8F",X"A6",X"49",X"74",X"75",X"AC",X"59",X"5D",X"67",X"9F",X"81",X"48",X"60",X"76",X"A8",
		X"3B",X"55",X"4E",X"BA",X"55",X"46",X"30",X"9B",X"86",X"3E",X"35",X"62",X"B4",X"51",X"5A",X"31",
		X"B0",X"74",X"77",X"42",X"74",X"A8",X"7C",X"7C",X"39",X"A8",X"90",X"A8",X"51",X"6A",X"B6",X"B3",
		X"9C",X"35",X"9C",X"A9",X"C9",X"63",X"5C",X"96",X"92",X"B2",X"3E",X"73",X"66",X"A8",X"8E",X"42",
		X"5D",X"50",X"BA",X"67",X"3A",X"2B",X"6F",X"B7",X"56",X"5F",X"2E",X"91",X"9B",X"72",X"78",X"37",
		X"A8",X"99",X"A7",X"6D",X"40",X"AF",X"B5",X"C9",X"5A",X"5B",X"A2",X"94",X"C0",X"4B",X"64",X"70",
		X"83",X"BD",X"4A",X"55",X"3B",X"81",X"B3",X"4C",X"54",X"31",X"87",X"B1",X"6B",X"87",X"35",X"84",
		X"AF",X"9D",X"A8",X"3A",X"7F",X"B5",X"B9",X"B0",X"3A",X"73",X"85",X"91",X"BD",X"45",X"5F",X"4D",
		X"74",X"C0",X"58",X"48",X"34",X"62",X"C1",X"75",X"82",X"57",X"45",X"B6",X"A0",X"C1",X"73",X"3F",
		X"9B",X"82",X"B6",X"96",X"3A",X"59",X"38",X"A2",X"AB",X"64",X"7F",X"38",X"72",X"BE",X"BB",X"C4",
		X"53",X"57",X"76",X"5A",X"C9",X"74",X"66",X"5F",X"42",X"86",X"43",X"38",X"32",X"33",X"33",X"32",
		X"33",X"33",X"34",X"33",X"35",X"34",X"36",X"35",X"37",X"36",X"39",X"37",X"39",X"38",X"3A",X"39",
		X"3B",X"3A",X"3B",X"3B",X"3B",X"3B",X"3C",X"3C",X"3D",X"3D",X"3D",X"3E",X"3F",X"3F",X"3F",X"40",
		X"40",X"41",X"41",X"42",X"42",X"42",X"42",X"43",X"43",X"44",X"44",X"45",X"45",X"46",X"46",X"47",
		X"47",X"48",X"48",X"49",X"49",X"49",X"4A",X"4A",X"4A",X"4A",X"4B",X"4B",X"4C",X"4C",X"4C",X"4D",
		X"4D",X"4D",X"4E",X"4E",X"4E",X"4F",X"4F",X"4F",X"50",X"50",X"50",X"51",X"50",X"51",X"51",X"51",
		X"51",X"52",X"52",X"53",X"53",X"53",X"54",X"54",X"55",X"55",X"56",X"56",X"56",X"57",X"57",X"57",
		X"58",X"58",X"58",X"58",X"58",X"59",X"59",X"59",X"5A",X"5A",X"5A",X"5A",X"5B",X"5B",X"5B",X"5B",
		X"5C",X"5C",X"5C",X"5C",X"5D",X"5D",X"5D",X"5D",X"5E",X"5E",X"5E",X"5E",X"5E",X"5E",X"5F",X"5F",
		X"5F",X"60",X"60",X"60",X"60",X"61",X"61",X"61",X"62",X"62",X"62",X"62",X"62",X"62",X"63",X"63",
		X"63",X"64",X"64",X"64",X"64",X"65",X"65",X"65",X"65",X"65",X"66",X"66",X"66",X"67",X"67",X"67",
		X"67",X"67",X"68",X"68",X"68",X"68",X"68",X"69",X"69",X"69",X"69",X"69",X"69",X"6A",X"6A",X"6A",
		X"6A",X"6A",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",
		X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"71",X"71",X"71",
		X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"73",X"73",X"73",X"73",X"73",X"73",X"73",
		X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"74",X"74",
		X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"75",X"75",X"75",X"75",X"76",X"76",
		X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",
		X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"78",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",
		X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",
		X"79",X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"80",X"81",X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"97",X"BE",X"B0",X"C0",X"BD",X"B5",X"C0",X"C1",X"D1",X"BF",X"D5",X"C5",X"C2",X"BC",X"BC",X"BE",
		X"A0",X"BC",X"B1",X"BB",X"BD",X"C2",X"CA",X"B7",X"D4",X"C6",X"BF",X"C6",X"B6",X"BE",X"AD",X"B9",
		X"B3",X"9D",X"B9",X"A6",X"A9",X"BA",X"AD",X"B7",X"B2",X"B5",X"BF",X"B2",X"C3",X"BD",X"B0",X"CE",
		X"BB",X"B8",X"D1",X"B2",X"B7",X"C6",X"AF",X"BB",X"BF",X"AB",X"B8",X"B7",X"AC",X"BA",X"B2",X"A9",
		X"B5",X"AE",X"AC",X"B6",X"AB",X"A8",X"B3",X"AA",X"A9",X"B5",X"AA",X"A5",X"B4",X"AD",X"A7",X"B9",
		X"B1",X"A1",X"B9",X"B9",X"A3",X"BE",X"C1",X"A0",X"B4",X"BD",X"A5",X"AB",X"B3",X"A3",X"9D",X"A8",
		X"A8",X"99",X"97",X"A6",X"93",X"84",X"A2",X"9E",X"88",X"98",X"A3",X"9C",X"9A",X"A6",X"B1",X"9F",
		X"9C",X"BD",X"B0",X"9A",X"A3",X"A5",X"9D",X"8A",X"91",X"A3",X"8F",X"80",X"98",X"9E",X"9C",X"94",
		X"A5",X"BA",X"A1",X"95",X"A2",X"A5",X"9B",X"84",X"89",X"9D",X"8F",X"8A",X"92",X"A6",X"AD",X"96",
		X"92",X"A4",X"A2",X"99",X"7D",X"88",X"99",X"95",X"90",X"8F",X"A4",X"B9",X"9B",X"8D",X"8A",X"95",
		X"9C",X"84",X"83",X"89",X"A5",X"A9",X"9A",X"8A",X"95",X"90",X"9C",X"79",X"87",X"87",X"AA",X"AB",
		X"96",X"86",X"85",X"91",X"95",X"8F",X"7D",X"8D",X"8D",X"B8",X"8D",X"9C",X"62",X"8B",X"82",X"A5",
		X"96",X"91",X"8B",X"84",X"9B",X"82",X"9C",X"6C",X"9E",X"76",X"B8",X"81",X"9C",X"6A",X"74",X"8F",
		X"89",X"CA",X"7B",X"A6",X"52",X"89",X"81",X"9B",X"B3",X"7E",X"9E",X"59",X"90",X"7F",X"9A",X"A8",
		X"7A",X"9B",X"5C",X"92",X"80",X"94",X"AB",X"76",X"9E",X"5E",X"87",X"89",X"86",X"B9",X"78",X"9B",
		X"6A",X"65",X"97",X"70",X"C3",X"90",X"87",X"8B",X"43",X"90",X"76",X"95",X"B3",X"74",X"9D",X"6E",
		X"6F",X"97",X"6C",X"9B",X"8D",X"78",X"A6",X"76",X"86",X"8E",X"52",X"8E",X"7A",X"84",X"C8",X"7B",
		X"93",X"84",X"50",X"90",X"76",X"78",X"A5",X"78",X"8F",X"AA",X"6C",X"93",X"76",X"42",X"92",X"76",
		X"85",X"B6",X"78",X"87",X"9C",X"6A",X"87",X"8D",X"4A",X"82",X"86",X"6C",X"B8",X"95",X"75",X"A3",
		X"82",X"68",X"9A",X"5F",X"4A",X"96",X"72",X"7E",X"AD",X"7B",X"77",X"AC",X"81",X"72",X"9E",X"57",
		X"54",X"93",X"6F",X"65",X"9C",X"81",X"71",X"C4",X"98",X"6C",X"97",X"87",X"61",X"89",X"84",X"39",
		X"72",X"8A",X"65",X"7E",X"9F",X"75",X"83",X"C6",X"8B",X"76",X"97",X"87",X"67",X"8A",X"82",X"41",
		X"6A",X"86",X"66",X"67",X"91",X"7A",X"70",X"A5",X"97",X"70",X"8C",X"AD",X"7F",X"7F",X"9E",X"7B",
		X"63",X"87",X"8E",X"45",X"5E",X"91",X"71",X"59",X"84",X"8A",X"5A",X"7D",X"A6",X"81",X"5E",X"A3",
		X"B9",X"6D",X"72",X"A0",X"91",X"62",X"87",X"9D",X"68",X"59",X"90",X"99",X"44",X"5C",X"95",X"8D",
		X"4F",X"6B",X"94",X"7A",X"5D",X"80",X"99",X"72",X"6B",X"93",X"9B",X"69",X"6D",X"A7",X"A2",X"69",
		X"6D",X"94",X"9C",X"63",X"71",X"7D",X"90",X"65",X"79",X"7D",X"7A",X"67",X"73",X"82",X"66",X"6D",
		X"70",X"8F",X"5B",X"63",X"6C",X"8B",X"64",X"62",X"73",X"88",X"73",X"6C",X"7A",X"81",X"76",X"71",
		X"85",X"87",X"7A",X"75",X"8E",X"8D",X"7B",X"6C",X"95",X"98",X"8B",X"64",X"92",X"9E",X"9B",X"60",
		X"7B",X"A6",X"A9",X"7B",X"5F",X"A6",X"AA",X"9F",X"4D",X"8D",X"AD",X"BB",X"6D",X"62",X"AB",X"B6",
		X"A3",X"45",X"8C",X"AF",X"C2",X"70",X"57",X"A8",X"B2",X"B0",X"46",X"7A",X"AC",X"BD",X"8C",X"45",
		X"9E",X"A6",X"BB",X"60",X"5B",X"A4",X"A8",X"AE",X"48",X"7C",X"9B",X"A7",X"92",X"41",X"8A",X"8E",
		X"AC",X"7B",X"4F",X"8E",X"81",X"A8",X"67",X"5B",X"82",X"7F",X"A4",X"63",X"66",X"71",X"79",X"98",
		X"61",X"5F",X"5E",X"79",X"94",X"69",X"57",X"50",X"71",X"8C",X"6C",X"4D",X"51",X"6D",X"8F",X"73",
		X"52",X"5E",X"61",X"8E",X"70",X"5D",X"70",X"5C",X"8E",X"78",X"6B",X"7C",X"55",X"84",X"81",X"7C",
		X"8F",X"58",X"7A",X"98",X"92",X"9D",X"5E",X"67",X"A2",X"92",X"AC",X"6F",X"5E",X"99",X"74",X"A6",
		X"83",X"51",X"89",X"61",X"95",X"A1",X"58",X"76",X"4E",X"71",X"AF",X"6B",X"55",X"42",X"4E",X"AD",
		X"85",X"5F",X"69",X"33",X"8C",X"9C",X"6B",X"94",X"47",X"5D",X"A7",X"85",X"AC",X"76",X"3A",X"84",
		X"A4",X"B9",X"B2",X"4B",X"60",X"98",X"85",X"BF",X"81",X"43",X"7B",X"60",X"8F",X"BB",X"5F",X"55",
		X"4C",X"48",X"AA",X"9D",X"54",X"57",X"39",X"64",X"B9",X"82",X"7C",X"76",X"37",X"82",X"AC",X"93",
		X"B1",X"68",X"44",X"94",X"AC",X"B3",X"B0",X"51",X"4F",X"8E",X"75",X"A7",X"A6",X"49",X"5C",X"5C",
		X"54",X"AD",X"95",X"4D",X"4C",X"3D",X"5A",X"B3",X"8B",X"6C",X"84",X"3E",X"63",X"A9",X"9D",X"AC",
		X"96",X"41",X"6D",X"97",X"7B",X"B3",X"8E",X"4A",X"57",X"4C",X"5D",X"B1",X"8E",X"65",X"80",X"46",
		X"5C",X"A1",X"AB",X"B2",X"A4",X"50",X"5E",X"79",X"58",X"9B",X"A5",X"5C",X"73",X"5D",X"4C",X"84",
		X"59",X"47",X"45",X"43",X"45",X"44",X"45",X"44",X"46",X"44",X"47",X"46",X"48",X"46",X"49",X"48",
		X"49",X"49",X"4B",X"4A",X"4B",X"4B",X"4C",X"4C",X"4D",X"4D",X"4D",X"4E",X"4E",X"4E",X"4E",X"4F",
		X"4F",X"50",X"50",X"51",X"51",X"52",X"52",X"53",X"53",X"53",X"54",X"54",X"54",X"55",X"55",X"56",
		X"56",X"56",X"57",X"57",X"58",X"58",X"58",X"59",X"59",X"5A",X"5A",X"5B",X"5B",X"5C",X"5C",X"5D",
		X"5D",X"5D",X"5E",X"5E",X"5E",X"5F",X"5F",X"5F",X"5F",X"60",X"60",X"61",X"61",X"61",X"61",X"62",
		X"62",X"62",X"63",X"63",X"63",X"64",X"64",X"64",X"64",X"65",X"65",X"65",X"65",X"66",X"66",X"66",
		X"66",X"66",X"66",X"67",X"67",X"67",X"68",X"68",X"68",X"68",X"69",X"69",X"69",X"6A",X"6A",X"6A",
		X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",
		X"6E",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"71",X"71",X"71",X"71",X"71",X"72",X"72",
		X"72",X"72",X"72",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",X"78",X"78",X"79",X"79",X"79",X"79",
		X"79",X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"80",X"81",X"81",X"80",X"80",
		X"80",X"81",X"80",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"80",X"80",X"81",X"7E",X"73",X"61",X"54",X"47",X"40",X"37",X"34",X"2D",X"3E",X"7B",X"95",
		X"96",X"98",X"96",X"96",X"94",X"94",X"93",X"8D",X"7B",X"6A",X"5C",X"51",X"4A",X"43",X"3F",X"3A",
		X"67",X"9C",X"A2",X"A4",X"A2",X"A1",X"9F",X"9E",X"9E",X"9B",X"90",X"7C",X"6C",X"5E",X"57",X"4E",
		X"4B",X"43",X"4E",X"8C",X"A9",X"A8",X"A9",X"A6",X"A6",X"A4",X"A3",X"A2",X"9E",X"8D",X"79",X"6B",
		X"5F",X"58",X"50",X"4E",X"45",X"68",X"A3",X"AD",X"AD",X"AB",X"AA",X"A8",X"A7",X"A6",X"A4",X"9B",
		X"86",X"76",X"69",X"5F",X"57",X"52",X"4D",X"4C",X"82",X"AD",X"AD",X"AE",X"AC",X"AB",X"A9",X"A7",
		X"A6",X"A3",X"95",X"81",X"73",X"65",X"5E",X"55",X"53",X"4A",X"59",X"97",X"AE",X"AD",X"AD",X"AA",
		X"A9",X"A6",X"A6",X"A5",X"9F",X"8E",X"7C",X"6D",X"62",X"5B",X"53",X"51",X"48",X"6B",X"A3",X"AC",
		X"AC",X"AA",X"A9",X"A7",X"A5",X"A4",X"A2",X"9A",X"87",X"76",X"68",X"5F",X"58",X"52",X"4E",X"4B",
		X"7C",X"A9",X"AA",X"AB",X"A8",X"A7",X"A4",X"A3",X"A1",X"9F",X"93",X"80",X"71",X"65",X"5D",X"55",
		X"51",X"4B",X"51",X"8A",X"A9",X"A8",X"A8",X"A5",X"A4",X"A2",X"A0",X"9E",X"9B",X"8C",X"79",X"6B",
		X"60",X"5A",X"53",X"51",X"49",X"57",X"92",X"A8",X"A7",X"A6",X"A3",X"A2",X"9F",X"9C",X"9A",X"95",
		X"86",X"74",X"67",X"5D",X"56",X"50",X"4F",X"47",X"5F",X"99",X"A6",X"A5",X"A3",X"A0",X"9D",X"9B",
		X"9A",X"98",X"92",X"82",X"71",X"65",X"5A",X"55",X"4E",X"4D",X"46",X"67",X"9E",X"A5",X"A4",X"A0",
		X"9E",X"9C",X"9A",X"99",X"97",X"90",X"7F",X"6F",X"62",X"59",X"53",X"4D",X"4C",X"46",X"6E",X"9F",
		X"A3",X"A2",X"9E",X"9D",X"9B",X"9A",X"98",X"97",X"8E",X"7D",X"6D",X"62",X"59",X"53",X"4D",X"4A",
		X"46",X"73",X"A0",X"A1",X"A1",X"9E",X"9D",X"9A",X"99",X"97",X"96",X"8D",X"7B",X"6C",X"61",X"58",
		X"53",X"4E",X"4B",X"48",X"77",X"A0",X"A1",X"A1",X"9D",X"9C",X"9A",X"99",X"97",X"96",X"8C",X"7B",
		X"6C",X"61",X"58",X"53",X"4E",X"4B",X"49",X"78",X"A0",X"A0",X"A0",X"9D",X"9C",X"99",X"99",X"97",
		X"95",X"8B",X"7B",X"6C",X"61",X"59",X"53",X"4E",X"4B",X"49",X"77",X"A0",X"A0",X"A0",X"9C",X"9C",
		X"99",X"99",X"97",X"96",X"8C",X"7B",X"6D",X"62",X"59",X"54",X"4E",X"4C",X"49",X"76",X"9F",X"A0",
		X"A0",X"9C",X"9C",X"99",X"98",X"96",X"96",X"8C",X"7C",X"6D",X"62",X"5A",X"55",X"4F",X"4D",X"49",
		X"72",X"9E",X"A0",X"A0",X"9C",X"9C",X"99",X"98",X"96",X"96",X"8D",X"7E",X"6F",X"64",X"5B",X"56",
		X"50",X"4E",X"49",X"6E",X"9C",X"A0",X"A0",X"9D",X"9C",X"99",X"98",X"97",X"96",X"8F",X"80",X"71",
		X"66",X"5D",X"57",X"51",X"50",X"49",X"66",X"99",X"A0",X"A0",X"9D",X"9C",X"99",X"99",X"97",X"96",
		X"91",X"82",X"73",X"68",X"5E",X"59",X"53",X"51",X"4A",X"5E",X"93",X"A0",X"A0",X"9E",X"9C",X"9A",
		X"99",X"97",X"96",X"92",X"85",X"76",X"6A",X"60",X"5A",X"54",X"52",X"4C",X"56",X"8B",X"A1",X"A0",
		X"9E",X"9C",X"9A",X"98",X"98",X"96",X"94",X"89",X"79",X"6C",X"63",X"5B",X"56",X"52",X"4F",X"50",
		X"80",X"A0",X"A0",X"9F",X"9C",X"9B",X"98",X"98",X"96",X"95",X"8C",X"7D",X"6F",X"65",X"5D",X"58",
		X"53",X"51",X"4D",X"72",X"9D",X"A0",X"A0",X"9C",X"9B",X"98",X"98",X"96",X"96",X"8F",X"81",X"72",
		X"68",X"5F",X"5A",X"55",X"53",X"4D",X"64",X"96",X"A0",X"A0",X"9D",X"9B",X"99",X"98",X"97",X"96",
		X"92",X"86",X"77",X"6C",X"62",X"5C",X"57",X"54",X"4F",X"57",X"89",X"A0",X"9F",X"9E",X"9B",X"9A",
		X"98",X"97",X"96",X"95",X"8A",X"7C",X"6F",X"66",X"5E",X"59",X"55",X"53",X"4F",X"77",X"9E",X"9F",
		X"9F",X"9B",X"9B",X"98",X"97",X"96",X"96",X"8F",X"81",X"73",X"69",X"61",X"5C",X"56",X"55",X"4F",
		X"63",X"95",X"A0",X"9F",X"9D",X"9B",X"99",X"97",X"96",X"95",X"93",X"87",X"79",X"6D",X"64",X"5E",
		X"59",X"56",X"52",X"54",X"82",X"A0",X"9F",X"9F",X"9B",X"9A",X"97",X"97",X"95",X"94",X"8D",X"7F",
		X"72",X"69",X"60",X"5C",X"56",X"55",X"4F",X"6A",X"99",X"A0",X"9F",X"9C",X"9B",X"98",X"97",X"95",
		X"94",X"91",X"85",X"77",X"6D",X"64",X"5E",X"59",X"56",X"53",X"57",X"86",X"A0",X"9F",X"9E",X"9B",
		X"99",X"96",X"96",X"94",X"94",X"8C",X"7E",X"71",X"69",X"61",X"5C",X"57",X"56",X"51",X"6C",X"99",
		X"9F",X"9F",X"9C",X"9A",X"97",X"96",X"95",X"94",X"91",X"85",X"77",X"6D",X"65",X"5F",X"5A",X"57",
		X"54",X"58",X"85",X"9F",X"9E",X"9D",X"9A",X"99",X"96",X"95",X"94",X"94",X"8C",X"7F",X"72",X"6A",
		X"61",X"5D",X"58",X"57",X"52",X"69",X"97",X"9F",X"9E",X"9B",X"9A",X"97",X"96",X"94",X"94",X"91",
		X"86",X"79",X"6E",X"66",X"60",X"5B",X"58",X"55",X"56",X"7F",X"9E",X"9E",X"9D",X"9A",X"99",X"96",
		X"95",X"93",X"94",X"8D",X"81",X"74",X"6B",X"63",X"5F",X"59",X"58",X"53",X"62",X"91",X"9F",X"9E",
		X"9C",X"99",X"98",X"95",X"95",X"93",X"92",X"89",X"7C",X"70",X"68",X"61",X"5D",X"59",X"58",X"53",
		X"73",X"9A",X"9E",X"9E",X"9A",X"99",X"96",X"95",X"94",X"93",X"8F",X"85",X"78",X"6E",X"66",X"60",
		X"5C",X"59",X"56",X"58",X"83",X"9E",X"9D",X"9D",X"99",X"98",X"96",X"95",X"93",X"93",X"8C",X"81",
		X"74",X"6B",X"64",X"5F",X"5A",X"59",X"54",X"62",X"8F",X"9E",X"9D",X"9C",X"99",X"97",X"95",X"94",
		X"92",X"92",X"89",X"7D",X"72",X"69",X"62",X"5F",X"5A",X"59",X"54",X"6D",X"97",X"9D",X"9D",X"9A",
		X"98",X"96",X"95",X"93",X"92",X"90",X"86",X"7A",X"6F",X"67",X"61",X"5E",X"5A",X"58",X"56",X"78",
		X"9B",X"9D",X"9C",X"99",X"98",X"95",X"94",X"93",X"92",X"8E",X"84",X"78",X"6E",X"66",X"61",X"5D",
		X"5A",X"57",X"5A",X"82",X"9D",X"9C",X"9C",X"99",X"98",X"94",X"94",X"92",X"92",X"8D",X"81",X"75",
		X"6C",X"65",X"61",X"5C",X"5B",X"57",X"5E",X"89",X"9D",X"9C",X"9B",X"98",X"97",X"94",X"94",X"92",
		X"91",X"8B",X"7F",X"74",X"6B",X"64",X"60",X"5C",X"5B",X"56",X"63",X"8F",X"9D",X"9C",X"9B",X"98",
		X"96",X"94",X"93",X"91",X"91",X"89",X"7E",X"73",X"6B",X"64",X"60",X"5C",X"5B",X"56",X"68",X"92",
		X"9D",X"9C",X"9A",X"98",X"96",X"94",X"93",X"91",X"90",X"88",X"7D",X"72",X"6A",X"64",X"60",X"5C",
		X"5C",X"56",X"6C",X"95",X"9C",X"9C",X"99",X"97",X"95",X"94",X"92",X"91",X"90",X"87",X"7C",X"71",
		X"6A",X"63",X"60",X"5C",X"5C",X"57",X"6F",X"96",X"9C",X"9B",X"99",X"97",X"95",X"94",X"92",X"91",
		X"8F",X"86",X"7B",X"71",X"6A",X"63",X"60",X"5D",X"5C",X"57",X"71",X"97",X"9B",X"9B",X"98",X"97",
		X"95",X"93",X"92",X"91",X"8F",X"86",X"7B",X"71",X"6A",X"64",X"60",X"5D",X"5C",X"58",X"71",X"97",
		X"9B",X"9B",X"98",X"96",X"94",X"93",X"92",X"90",X"8F",X"86",X"7B",X"71",X"6A",X"64",X"61",X"5D",
		X"5C",X"58",X"71",X"96",X"9B",X"9A",X"98",X"96",X"94",X"93",X"92",X"90",X"8F",X"87",X"7B",X"71",
		X"6B",X"64",X"61",X"5D",X"5D",X"59",X"6F",X"95",X"9B",X"9A",X"98",X"96",X"94",X"93",X"91",X"90",
		X"8F",X"87",X"7C",X"72",X"6B",X"65",X"62",X"5E",X"5D",X"59",X"6C",X"93",X"9B",X"9A",X"98",X"96",
		X"94",X"93",X"91",X"90",X"8F",X"88",X"7D",X"73",X"6C",X"66",X"62",X"5E",X"5E",X"5A",X"68",X"8F",
		X"9B",X"9A",X"98",X"96",X"95",X"93",X"92",X"90",X"8F",X"89",X"7F",X"74",X"6D",X"66",X"63",X"5F",
		X"5E",X"5A",X"63",X"8A",X"9B",X"99",X"98",X"96",X"95",X"92",X"92",X"90",X"90",X"8A",X"80",X"76",
		X"6E",X"68",X"64",X"60",X"5F",X"5C",X"5F",X"84",X"9A",X"99",X"99",X"96",X"95",X"93",X"92",X"90",
		X"90",X"8C",X"82",X"78",X"70",X"69",X"64",X"61",X"5F",X"5E",X"5C",X"7B",X"99",X"99",X"99",X"96",
		X"95",X"93",X"92",X"90",X"8F",X"8D",X"84",X"7A",X"71",X"6B",X"65",X"62",X"5F",X"5F",X"5B",X"71",
		X"94",X"9A",X"99",X"97",X"95",X"94",X"92",X"90",X"8F",X"8E",X"87",X"7D",X"73",X"6D",X"67",X"64",
		X"60",X"5F",X"5B",X"68",X"8D",X"9A",X"99",X"97",X"95",X"94",X"92",X"91",X"8F",X"8F",X"8A",X"80",
		X"76",X"6F",X"68",X"65",X"61",X"60",X"5D",X"60",X"83",X"99",X"98",X"98",X"96",X"95",X"92",X"91",
		X"8F",X"8F",X"8C",X"83",X"79",X"71",X"6B",X"65",X"63",X"60",X"5F",X"5D",X"76",X"96",X"99",X"98",
		X"96",X"95",X"93",X"91",X"90",X"8F",X"8D",X"86",X"7C",X"73",X"6D",X"67",X"64",X"61",X"60",X"5D",
		X"6A",X"8D",X"99",X"98",X"97",X"95",X"93",X"91",X"91",X"8F",X"8E",X"89",X"80",X"76",X"6F",X"69",
		X"66",X"62",X"60",X"5F",X"61",X"82",X"98",X"97",X"98",X"95",X"94",X"92",X"91",X"8F",X"8E",X"8B",
		X"83",X"79",X"71",X"6B",X"66",X"64",X"61",X"60",X"5E",X"77",X"95",X"98",X"98",X"95",X"94",X"92",
		X"91",X"8F",X"8E",X"8D",X"85",X"7B",X"73",X"6D",X"67",X"64",X"61",X"61",X"5D",X"72",X"93",X"98",
		X"97",X"95",X"94",X"92",X"91",X"8F",X"8E",X"8D",X"86",X"7C",X"73",X"6D",X"67",X"65",X"62",X"61",
		X"5E",X"72",X"93",X"97",X"96",X"95",X"93",X"92",X"90",X"8F",X"8E",X"8C",X"85",X"7B",X"73",X"6C",
		X"68",X"65",X"62",X"61",X"5F",X"78",X"95",X"97",X"96",X"94",X"93",X"91",X"90",X"8E",X"8D",X"8B",
		X"83",X"79",X"72",X"6B",X"67",X"64",X"63",X"60",X"63",X"83",X"97",X"96",X"95",X"93",X"92",X"90",
		X"8F",X"8D",X"8D",X"88",X"7F",X"76",X"6F",X"69",X"67",X"64",X"62",X"5F",X"6F",X"90",X"96",X"96",
		X"94",X"92",X"91",X"8F",X"8E",X"8E",X"8B",X"84",X"7A",X"72",X"6C",X"68",X"66",X"63",X"61",X"64",
		X"84",X"96",X"95",X"95",X"93",X"91",X"90",X"8F",X"8D",X"8C",X"86",X"7D",X"75",X"6F",X"6A",X"67",
		X"64",X"63",X"61",X"7A",X"94",X"95",X"95",X"93",X"92",X"90",X"8F",X"8D",X"8D",X"88",X"7F",X"77",
		X"70",X"6B",X"68",X"64",X"63",X"60",X"74",X"92",X"96",X"95",X"93",X"91",X"90",X"8F",X"8D",X"8C",
		X"89",X"80",X"77",X"71",X"6B",X"68",X"65",X"64",X"60",X"72",X"90",X"96",X"95",X"93",X"91",X"90",
		X"8F",X"8D",X"8C",X"89",X"80",X"77",X"71",X"6B",X"68",X"65",X"64",X"61",X"75",X"91",X"95",X"95",
		X"92",X"91",X"90",X"8E",X"8D",X"8C",X"88",X"7F",X"76",X"70",X"6B",X"68",X"65",X"64",X"62",X"7B",
		X"93",X"94",X"94",X"92",X"91",X"8F",X"8E",X"8D",X"8B",X"86",X"7D",X"75",X"6E",X"6B",X"67",X"65",
		X"63",X"66",X"84",X"94",X"94",X"94",X"91",X"90",X"8E",X"8D",X"8C",X"8A",X"83",X"7A",X"73",X"6D",
		X"6A",X"66",X"66",X"62",X"70",X"8E",X"94",X"93",X"92",X"90",X"8F",X"8E",X"8D",X"8B",X"88",X"7F",
		X"77",X"70",X"6B",X"68",X"66",X"64",X"65",X"81",X"94",X"93",X"93",X"90",X"90",X"8E",X"8D",X"8C",
		X"8A",X"83",X"7A",X"73",X"6D",X"6A",X"67",X"65",X"62",X"74",X"8F",X"94",X"93",X"92",X"90",X"8F",
		X"8D",X"8C",X"8B",X"86",X"7D",X"75",X"6F",X"6C",X"68",X"66",X"63",X"6C",X"89",X"93",X"93",X"92",
		X"90",X"8F",X"8D",X"8C",X"8B",X"87",X"7F",X"77",X"71",X"6C",X"68",X"67",X"64",X"68",X"83",X"93",
		X"93",X"92",X"90",X"8F",X"8D",X"8C",X"8B",X"88",X"80",X"78",X"72",X"6D",X"69",X"67",X"65",X"66",
		X"80",X"93",X"92",X"92",X"90",X"8F",X"8D",X"8C",X"8B",X"88",X"81",X"79",X"72",X"6D",X"6A",X"68",
		X"65",X"66",X"81",X"92",X"92",X"92",X"8F",X"8F",X"8D",X"8C",X"8B",X"88",X"80",X"78",X"72",X"6D",
		X"6A",X"68",X"65",X"68",X"83",X"93",X"92",X"91",X"8F",X"8E",X"8D",X"8C",X"8B",X"88",X"7F",X"77",
		X"71",X"6D",X"69",X"67",X"64",X"6C",X"88",X"92",X"92",X"91",X"8F",X"8E",X"8C",X"8C",X"8A",X"85",
		X"7D",X"76",X"70",X"6C",X"68",X"68",X"64",X"73",X"8D",X"92",X"91",X"90",X"8F",X"8D",X"8C",X"8B",
		X"8A",X"83",X"7A",X"74",X"6F",X"6B",X"68",X"67",X"66",X"7E",X"91",X"91",X"91",X"8F",X"8E",X"8C",
		X"8C",X"8B",X"87",X"7F",X"78",X"71",X"6E",X"6A",X"69",X"65",X"6E",X"8A",X"91",X"91",X"90",X"8E",
		X"8D",X"8C",X"8B",X"89",X"83",X"7B",X"75",X"6F",X"6C",X"69",X"67",X"67",X"7E",X"91",X"91",X"91",
		X"8F",X"8D",X"8C",X"8B",X"8A",X"87",X"7E",X"77",X"71",X"6E",X"6A",X"69",X"65",X"74",X"8D",X"91",
		X"90",X"8F",X"8E",X"8C",X"8B",X"8A",X"88",X"81",X"79",X"73",X"6F",X"6B",X"69",X"66",X"6D",X"88",
		X"91",X"90",X"8F",X"8E",X"8C",X"8B",X"8B",X"89",X"83",X"7B",X"75",X"6F",X"6C",X"69",X"67",X"6A",
		X"84",X"90",X"90",X"90",X"8D",X"8D",X"8C",X"8B",X"89",X"84",X"7C",X"75",X"70",X"6D",X"6A",X"68",
		X"69",X"81",X"90",X"90",X"90",X"8D",X"8D",X"8C",X"8B",X"89",X"84",X"7C",X"76",X"70",X"6D",X"6A",
		X"68",X"69",X"80",X"90",X"90",X"90",X"8E",X"8D",X"8B",X"8B",X"89",X"84",X"7C",X"76",X"71",X"6D",
		X"6B",X"69",X"69",X"80",X"90",X"90",X"8F",X"8E",X"8D",X"8B",X"8B",X"89",X"83",X"7C",X"75",X"71",
		X"6D",X"6B",X"68",X"6B",X"83",X"90",X"90",X"8F",X"8D",X"8C",X"8B",X"8A",X"88",X"82",X"7B",X"74",
		X"70",X"6C",X"6B",X"68",X"6E",X"87",X"90",X"8F",X"8F",X"8D",X"8C",X"8B",X"8A",X"87",X"80",X"79",
		X"74",X"6F",X"6C",X"6A",X"67",X"74",X"8B",X"90",X"8F",X"8E",X"8C",X"8C",X"8A",X"8A",X"86",X"7E",
		X"77",X"72",X"6E",X"6C",X"69",X"69",X"7D",X"8F",X"8F",X"8F",X"8D",X"8C",X"8B",X"8A",X"89",X"83",
		X"7C",X"75",X"71",X"6D",X"6B",X"68",X"6F",X"87",X"90",X"8E",X"8E",X"8C",X"8C",X"8A",X"8A",X"86",
		X"80",X"79",X"73",X"6F",X"6C",X"6A",X"68",X"7B",X"8E",X"8F",X"8F",X"8D",X"8C",X"8B",X"8A",X"89",
		X"83",X"7C",X"76",X"71",X"6D",X"6C",X"68",X"70",X"88",X"8F",X"8E",X"8E",X"8C",X"8B",X"8A",X"89",
		X"85",X"7F",X"78",X"73",X"6F",X"6C",X"6A",X"6B",X"7F",X"8E",X"8E",X"8E",X"8C",X"8C",X"8A",X"8A",
		X"87",X"81",X"7B",X"75",X"71",X"6D",X"6B",X"69",X"77",X"8B",X"8E",X"8E",X"8D",X"8C",X"8B",X"8A",
		X"89",X"84",X"7D",X"77",X"72",X"6E",X"6D",X"69",X"6F",X"86",X"8F",X"8E",X"8D",X"8C",X"8B",X"8A",
		X"89",X"86",X"80",X"79",X"74",X"70",X"6D",X"6B",X"6A",X"7D",X"8E",X"8E",X"8E",X"8C",X"8B",X"8A",
		X"89",X"88",X"82",X"7B",X"75",X"71",X"6E",X"6C",X"69",X"73",X"8A",X"8E",X"8D",X"8D",X"8B",X"8B",
		X"89",X"89",X"85",X"7E",X"78",X"73",X"6F",X"6D",X"6A",X"6C",X"80",X"8E",X"8E",X"8D",X"8C",X"8B",
		X"8A",X"89",X"87",X"81",X"7A",X"75",X"71",X"6E",X"6C",X"69",X"75",X"8A",X"8E",X"8D",X"8C",X"8B",
		X"8B",X"89",X"89",X"85",X"7E",X"78",X"73",X"6F",X"6D",X"6B",X"6C",X"81",X"8E",X"8D",X"8D",X"8C",
		X"8B",X"8A",X"89",X"87",X"82",X"7B",X"75",X"71",X"6E",X"6D",X"69",X"74",X"89",X"8E",X"8D",X"8C",
		X"8B",X"8A",X"89",X"89",X"85",X"7F",X"78",X"74",X"70",X"6E",X"6C",X"6B",X"7E",X"8D",X"8D",X"8D",
		X"8C",X"8B",X"8A",X"89",X"88",X"82",X"7C",X"76",X"72",X"6E",X"6D",X"6A",X"71",X"86",X"8E",X"8D",
		X"8D",X"8B",X"8B",X"89",X"89",X"86",X"80",X"7A",X"74",X"71",X"6E",X"6D",X"6A",X"79",X"8B",X"8E",
		X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"84",X"7E",X"78",X"73",X"70",X"6E",X"6B",X"6D",X"81",X"8D",
		X"8D",X"8D",X"8B",X"8A",X"89",X"89",X"87",X"82",X"7C",X"76",X"72",X"6F",X"6E",X"6B",X"72",X"87",
		X"8E",X"8D",X"8D",X"8B",X"8A",X"89",X"89",X"86",X"80",X"7A",X"75",X"72",X"6F",X"6D",X"6B",X"77",
		X"8B",X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"85",X"7F",X"79",X"74",X"71",X"6F",X"6D",X"6C",
		X"7D",X"8C",X"8D",X"8D",X"8B",X"8A",X"89",X"89",X"88",X"84",X"7D",X"78",X"73",X"70",X"6E",X"6C",
		X"6E",X"81",X"8D",X"8D",X"8D",X"8B",X"8A",X"89",X"89",X"87",X"83",X"7C",X"77",X"73",X"70",X"6E",
		X"6C",X"70",X"85",X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"87",X"81",X"7B",X"76",X"72",X"6F",
		X"6E",X"6B",X"72",X"87",X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"86",X"81",X"7B",X"75",X"72",
		X"6F",X"6E",X"6B",X"74",X"88",X"8D",X"8D",X"8B",X"8A",X"8A",X"88",X"88",X"86",X"80",X"7A",X"75",
		X"72",X"6F",X"6E",X"6B",X"75",X"89",X"8D",X"8D",X"8B",X"8A",X"89",X"88",X"88",X"86",X"80",X"7A",
		X"75",X"72",X"6F",X"6E",X"6C",X"76",X"89",X"8D",X"8D",X"8B",X"8A",X"89",X"88",X"88",X"86",X"80",
		X"7A",X"75",X"72",X"6F",X"6E",X"6C",X"76",X"89",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"88",X"86",
		X"80",X"7A",X"75",X"72",X"6F",X"6F",X"6C",X"75",X"88",X"8C",X"8C",X"8B",X"8A",X"89",X"88",X"88",
		X"86",X"80",X"7B",X"76",X"73",X"70",X"6F",X"6C",X"74",X"88",X"8C",X"8C",X"8B",X"8A",X"89",X"88",
		X"87",X"86",X"81",X"7B",X"76",X"73",X"70",X"6F",X"6D",X"73",X"86",X"8C",X"8C",X"8B",X"8A",X"89",
		X"88",X"87",X"86",X"82",X"7C",X"77",X"73",X"71",X"6F",X"6D",X"72",X"84",X"8C",X"8C",X"8B",X"8A",
		X"89",X"88",X"87",X"87",X"82",X"7C",X"77",X"74",X"71",X"70",X"6E",X"70",X"83",X"8C",X"8C",X"8B",
		X"8A",X"89",X"88",X"88",X"87",X"82",X"7C",X"78",X"74",X"71",X"70",X"6E",X"6F",X"81",X"8C",X"8C",
		X"8B",X"8A",X"89",X"88",X"88",X"87",X"83",X"7D",X"78",X"74",X"72",X"70",X"6E",X"6F",X"81",X"8C",
		X"8C",X"8B",X"8A",X"89",X"88",X"88",X"87",X"82",X"7D",X"78",X"74",X"72",X"70",X"6E",X"70",X"82",
		X"8C",X"8C",X"8B",X"8A",X"89",X"88",X"88",X"86",X"82",X"7C",X"77",X"74",X"71",X"70",X"6E",X"71",
		X"84",X"8C",X"8B",X"8B",X"8A",X"89",X"88",X"87",X"86",X"81",X"7B",X"76",X"73",X"71",X"70",X"6E",
		X"75",X"87",X"8C",X"8B",X"8B",X"89",X"89",X"88",X"87",X"85",X"7F",X"7A",X"75",X"73",X"71",X"6F",
		X"6E",X"7B",X"8A",X"8C",X"8B",X"8A",X"89",X"89",X"87",X"87",X"83",X"7D",X"78",X"74",X"72",X"70",
		X"6E",X"71",X"83",X"8B",X"8B",X"8B",X"89",X"89",X"88",X"87",X"85",X"81",X"7B",X"76",X"74",X"71",
		X"70",X"6E",X"79",X"89",X"8B",X"8B",X"8A",X"89",X"88",X"88",X"87",X"83",X"7E",X"79",X"75",X"72",
		X"71",X"6F",X"72",X"82",X"8B",X"8B",X"8B",X"89",X"89",X"88",X"87",X"85",X"80",X"7B",X"77",X"74",
		X"71",X"70",X"6F",X"7B",X"89",X"8B",X"8B",X"8A",X"89",X"88",X"87",X"86",X"82",X"7C",X"78",X"75",
		X"72",X"71",X"6F",X"75",X"86",X"8B",X"8A",X"8A",X"89",X"88",X"87",X"87",X"83",X"7E",X"79",X"76",
		X"73",X"71",X"6F",X"72",X"82",X"8B",X"8A",X"8A",X"89",X"88",X"87",X"87",X"84",X"7F",X"7A",X"76",
		X"74",X"72",X"70",X"71",X"7F",X"8A",X"8A",X"8A",X"89",X"88",X"87",X"87",X"85",X"80",X"7B",X"77",
		X"74",X"72",X"70",X"70",X"7D",X"8A",X"8A",X"8A",X"89",X"88",X"87",X"87",X"85",X"81",X"7B",X"77",
		X"74",X"72",X"71",X"70",X"7C",X"89",X"8A",X"8A",X"89",X"88",X"87",X"87",X"85",X"81",X"7C",X"77",
		X"75",X"72",X"71",X"70",X"7C",X"89",X"8A",X"8A",X"88",X"88",X"87",X"87",X"85",X"80",X"7B",X"77",
		X"74",X"72",X"71",X"71",X"7E",X"89",X"8A",X"89",X"88",X"88",X"87",X"87",X"84",X"80",X"7B",X"77",
		X"74",X"72",X"71",X"71",X"80",X"8A",X"8A",X"89",X"88",X"88",X"87",X"86",X"84",X"7F",X"7A",X"77",
		X"74",X"72",X"70",X"73",X"83",X"8A",X"8A",X"89",X"88",X"88",X"87",X"86",X"83",X"7E",X"7A",X"76",
		X"73",X"72",X"70",X"76",X"85",X"8A",X"89",X"89",X"88",X"87",X"86",X"86",X"82",X"7D",X"78",X"76",
		X"73",X"72",X"70",X"7B",X"88",X"89",X"89",X"88",X"88",X"87",X"86",X"84",X"80",X"7B",X"77",X"75",
		X"73",X"71",X"73",X"81",X"89",X"89",X"89",X"88",X"87",X"87",X"86",X"83",X"7E",X"7A",X"77",X"74",
		X"73",X"70",X"78",X"86",X"89",X"89",X"88",X"87",X"87",X"86",X"85",X"81",X"7C",X"78",X"75",X"73",
		X"72",X"72",X"7F",X"89",X"89",X"89",X"87",X"87",X"86",X"86",X"83",X"7E",X"7A",X"77",X"74",X"73",
		X"70",X"78",X"86",X"89",X"89",X"88",X"87",X"87",X"86",X"85",X"81",X"7C",X"78",X"75",X"73",X"71",
		X"73",X"81",X"89",X"89",X"89",X"87",X"87",X"86",X"85",X"82",X"7E",X"79",X"77",X"74",X"73",X"71",
		X"7B",X"88",X"89",X"89",X"88",X"87",X"86",X"86",X"83",X"7F",X"7B",X"78",X"75",X"73",X"71",X"77",
		X"85",X"89",X"89",X"88",X"87",X"86",X"86",X"84",X"81",X"7C",X"78",X"76",X"74",X"72",X"74",X"82",
		X"89",X"89",X"88",X"87",X"86",X"86",X"85",X"81",X"7D",X"79",X"76",X"74",X"72",X"73",X"80",X"88",
		X"88",X"88",X"87",X"87",X"86",X"85",X"82",X"7E",X"79",X"77",X"74",X"73",X"72",X"7E",X"88",X"88",
		X"88",X"87",X"87",X"86",X"86",X"83",X"7E",X"7A",X"77",X"74",X"73",X"71",X"7D",X"88",X"88",X"88",
		X"87",X"87",X"86",X"85",X"83",X"7E",X"7A",X"77",X"75",X"73",X"72",X"7C",X"88",X"88",X"88",X"87",
		X"87",X"86",X"85",X"83",X"7F",X"7A",X"77",X"75",X"73",X"72",X"7C",X"87",X"88",X"88",X"87",X"87",
		X"85",X"85",X"82",X"7E",X"7A",X"77",X"75",X"74",X"72",X"7D",X"87",X"88",X"88",X"87",X"87",X"85",
		X"85",X"82",X"7E",X"7A",X"77",X"75",X"73",X"73",X"7F",X"88",X"88",X"87",X"86",X"86",X"85",X"84",
		X"82",X"7D",X"7A",X"76",X"75",X"73",X"74",X"80",X"88",X"88",X"88",X"87",X"86",X"85",X"84",X"81",
		X"7C",X"79",X"76",X"74",X"72",X"75",X"82",X"88",X"88",X"87",X"87",X"86",X"85",X"84",X"80",X"7B",
		X"79",X"76",X"74",X"72",X"78",X"85",X"88",X"88",X"87",X"86",X"85",X"85",X"83",X"7F",X"7B",X"78",
		X"75",X"74",X"72",X"7B",X"87",X"88",X"88",X"87",X"86",X"85",X"85",X"83",X"7E",X"7A",X"77",X"75",
		X"74",X"73",X"7D",X"87",X"88",X"87",X"87",X"86",X"85",X"85",X"82",X"7E",X"7A",X"77",X"75",X"73",
		X"73",X"7F",X"88",X"87",X"87",X"86",X"86",X"85",X"84",X"81",X"7D",X"7A",X"77",X"75",X"74",X"75",
		X"80",X"88",X"88",X"87",X"86",X"85",X"85",X"84",X"81",X"7D",X"7A",X"77",X"75",X"73",X"75",X"82",
		X"88",X"88",X"87",X"87",X"86",X"85",X"84",X"80",X"7C",X"79",X"77",X"75",X"73",X"75",X"82",X"87",
		X"87",X"87",X"87",X"86",X"86",X"85",X"81",X"7C",X"79",X"77",X"75",X"73",X"75",X"82",X"87",X"87",
		X"87",X"86",X"86",X"85",X"84",X"81",X"7D",X"7A",X"78",X"76",X"74",X"76",X"82",X"87",X"87",X"86",
		X"86",X"85",X"85",X"84",X"80",X"7D",X"7B",X"78",X"77",X"75",X"77",X"82",X"87",X"87",X"87",X"86",
		X"85",X"83",X"83",X"82",X"88",X"93",X"97",X"96",X"95",X"92",X"86",X"7E",X"7D",X"7C",X"7C",X"7D",
		X"7D",X"7E",X"88",X"90",X"91",X"90",X"8F",X"8E",X"8D",X"81",X"76",X"76",X"76",X"77",X"77",X"78",
		X"79",X"83",X"8C",X"8E",X"8D",X"8B",X"8A",X"8A",X"80",X"73",X"72",X"72",X"73",X"73",X"75",X"75",
		X"7D",X"89",X"8C",X"8B",X"8A",X"89",X"89",X"81",X"73",X"70",X"70",X"71",X"72",X"72",X"73",X"79",
		X"85",X"8A",X"8A",X"89",X"88",X"88",X"84",X"76",X"70",X"70",X"70",X"71",X"72",X"72",X"75",X"81",
		X"89",X"8A",X"89",X"88",X"88",X"87",X"7B",X"70",X"70",X"70",X"72",X"72",X"73",X"73",X"7D",X"88",
		X"8A",X"8A",X"89",X"88",X"88",X"81",X"73",X"70",X"70",X"71",X"72",X"73",X"73",X"78",X"84",X"8B",
		X"8B",X"8A",X"88",X"88",X"86",X"79",X"70",X"71",X"71",X"72",X"73",X"73",X"74",X"7F",X"8A",X"8C",
		X"8B",X"8A",X"89",X"89",X"81",X"74",X"71",X"72",X"73",X"73",X"74",X"75",X"79",X"85",X"8B",X"8B",
		X"8B",X"8A",X"89",X"88",X"7B",X"72",X"72",X"72",X"74",X"74",X"76",X"76",X"7E",X"89",X"8D",X"8C",
		X"8B",X"8A",X"89",X"84",X"76",X"72",X"72",X"73",X"74",X"75",X"76",X"78",X"84",X"8C",X"8D",X"8C",
		X"8B",X"8A",X"8A",X"80",X"74",X"73",X"73",X"74",X"75",X"76",X"77",X"7C",X"88",X"8D",X"8D",X"8D",
		X"8C",X"8B",X"89",X"7C",X"73",X"73",X"73",X"75",X"76",X"77",X"77",X"7F",X"8B",X"8E",X"8E",X"8D",
		X"8C",X"8B",X"87",X"79",X"73",X"74",X"75",X"76",X"76",X"77",X"78",X"82",X"8C",X"8F",X"8E",X"8D",
		X"8B",X"8B",X"85",X"77",X"73",X"74",X"75",X"76",X"77",X"77",X"79",X"84",X"8D",X"8F",X"8D",X"8C",
		X"8B",X"8B",X"83",X"76",X"73",X"74",X"75",X"76",X"77",X"78",X"7A",X"85",X"8E",X"8F",X"8D",X"8C",
		X"8B",X"8B",X"82",X"75",X"74",X"74",X"75",X"76",X"77",X"77",X"7B",X"86",X"8E",X"8F",X"8D",X"8C",
		X"8B",X"8A",X"81",X"75",X"74",X"74",X"75",X"76",X"77",X"77",X"7B",X"86",X"8E",X"8E",X"8D",X"8C",
		X"8B",X"8A",X"81",X"75",X"74",X"74",X"75",X"76",X"77",X"77",X"7A",X"86",X"8E",X"8E",X"8D",X"8C",
		X"8B",X"8B",X"82",X"75",X"73",X"74",X"75",X"76",X"77",X"77",X"7A",X"84",X"8D",X"8F",X"8D",X"8C",
		X"8B",X"8B",X"84",X"76",X"73",X"74",X"75",X"76",X"76",X"77",X"79",X"82",X"8C",X"8F",X"8E",X"8D",
		X"8B",X"8B",X"86",X"78",X"73",X"74",X"75",X"76",X"76",X"77",X"78",X"7F",X"8B",X"8F",X"8E",X"8D",
		X"8B",X"8B",X"88",X"7B",X"73",X"73",X"74",X"75",X"76",X"77",X"77",X"7C",X"88",X"8E",X"8E",X"8D",
		X"8C",X"8B",X"8A",X"7F",X"74",X"73",X"74",X"75",X"76",X"77",X"77",X"7A",X"84",X"8D",X"8E",X"8D",
		X"8C",X"8B",X"8B",X"84",X"76",X"73",X"73",X"74",X"76",X"76",X"77",X"78",X"80",X"8B",X"8E",X"8E",
		X"8D",X"8B",X"8B",X"88",X"7B",X"73",X"73",X"74",X"75",X"76",X"77",X"77",X"7B",X"87",X"8D",X"8E",
		X"8D",X"8C",X"8A",X"8A",X"82",X"75",X"73",X"74",X"75",X"76",X"76",X"77",X"78",X"81",X"8B",X"8E",
		X"8D",X"8C",X"8B",X"8A",X"88",X"7B",X"73",X"73",X"74",X"75",X"76",X"77",X"77",X"7B",X"86",X"8D",
		X"8E",X"8D",X"8C",X"8A",X"8A",X"83",X"76",X"73",X"74",X"75",X"75",X"76",X"77",X"78",X"7F",X"8A",
		X"8E",X"8D",X"8C",X"8B",X"8A",X"89",X"7D",X"73",X"73",X"74",X"75",X"76",X"77",X"77",X"79",X"83",
		X"8C",X"8E",X"8D",X"8C",X"8B",X"8A",X"87",X"79",X"73",X"73",X"74",X"75",X"76",X"77",X"77",X"7B",
		X"86",X"8D",X"8E",X"8D",X"8C",X"8A",X"8A",X"84",X"76",X"73",X"74",X"74",X"75",X"76",X"77",X"77",
		X"7D",X"88",X"8D",X"8E",X"8C",X"8B",X"8A",X"8A",X"81",X"75",X"73",X"74",X"75",X"75",X"76",X"77",
		X"78",X"7F",X"8A",X"8E",X"8D",X"8C",X"8B",X"8A",X"8A",X"7F",X"74",X"73",X"74",X"75",X"75",X"76",
		X"77",X"78",X"80",X"8A",X"8E",X"8D",X"8C",X"8B",X"8A",X"89",X"7E",X"73",X"73",X"74",X"75",X"75",
		X"76",X"77",X"79",X"81",X"8B",X"8E",X"8D",X"8C",X"8B",X"8A",X"89",X"7D",X"73",X"73",X"74",X"75",
		X"76",X"77",X"77",X"79",X"81",X"8B",X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"7D",X"73",X"73",X"74",
		X"75",X"75",X"77",X"77",X"79",X"80",X"8A",X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"7E",X"74",X"73",
		X"74",X"75",X"75",X"77",X"77",X"78",X"7F",X"8A",X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"80",X"74",
		X"73",X"74",X"75",X"75",X"77",X"77",X"78",X"7D",X"88",X"8D",X"8D",X"8C",X"8C",X"8A",X"8A",X"83",
		X"76",X"73",X"74",X"75",X"75",X"76",X"77",X"78",X"7B",X"86",X"8D",X"8D",X"8C",X"8C",X"8B",X"8A",
		X"86",X"78",X"73",X"73",X"74",X"75",X"76",X"77",X"77",X"7A",X"82",X"8B",X"8D",X"8D",X"8C",X"8B",
		X"8A",X"88",X"7D",X"74",X"73",X"74",X"75",X"76",X"77",X"77",X"78",X"7E",X"89",X"8D",X"8D",X"8C",
		X"8B",X"8A",X"8A",X"82",X"76",X"73",X"74",X"75",X"75",X"77",X"77",X"78",X"7B",X"85",X"8C",X"8D",
		X"8D",X"8C",X"8A",X"8A",X"87",X"7A",X"73",X"73",X"74",X"75",X"76",X"77",X"77",X"79",X"7F",X"8A",
		X"8D",X"8D",X"8C",X"8B",X"8A",X"8A",X"81",X"75",X"73",X"74",X"75",X"75",X"77",X"77",X"78",X"7B",
		X"85",X"8C",X"8D",X"8D",X"8C",X"8A",X"8A",X"87",X"7B",X"73",X"73",X"74",X"75",X"76",X"77",X"77",
		X"78",X"7F",X"88",X"8D",X"8D",X"8C",X"8B",X"8A",X"8A",X"83",X"76",X"73",X"74",X"75",X"76",X"76",
		X"77",X"78",X"7A",X"82",X"8B",X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"7E",X"74",X"73",X"74",X"75",
		X"76",X"77",X"77",X"78",X"7C",X"85",X"8C",X"8D",X"8C",X"8C",X"8A",X"8A",X"87",X"7B",X"73",X"74",
		X"74",X"75",X"76",X"77",X"78",X"78",X"7E",X"87",X"8C",X"8D",X"8C",X"8C",X"8A",X"8A",X"85",X"78",
		X"73",X"74",X"75",X"76",X"76",X"77",X"78",X"79",X"7F",X"89",X"8D",X"8D",X"8C",X"8B",X"8A",X"8A",
		X"84",X"77",X"73",X"74",X"75",X"76",X"77",X"77",X"78",X"79",X"80",X"89",X"8D",X"8D",X"8C",X"8B",
		X"8A",X"89",X"83",X"76",X"73",X"74",X"75",X"76",X"77",X"77",X"78",X"79",X"80",X"8A",X"8D",X"8D",
		X"8C",X"8B",X"8A",X"89",X"83",X"76",X"73",X"74",X"75",X"76",X"77",X"78",X"78",X"79",X"80",X"89",
		X"8D",X"8D",X"8C",X"8B",X"8A",X"89",X"83",X"76",X"73",X"74",X"75",X"76",X"77",X"78",X"78",X"79",
		X"80",X"89",X"8D",X"8D",X"8C",X"8B",X"8A",X"8A",X"84",X"77",X"73",X"74",X"75",X"76",X"76",X"78",
		X"78",X"79",X"7F",X"88",X"8C",X"8D",X"8C",X"8B",X"8A",X"8A",X"86",X"79",X"73",X"74",X"74",X"75",
		X"76",X"77",X"78",X"79",X"7D",X"86",X"8C",X"8D",X"8C",X"8B",X"8A",X"89",X"87",X"7B",X"73",X"74",
		X"74",X"75",X"76",X"77",X"78",X"78",X"7B",X"84",X"8B",X"8D",X"8D",X"8C",X"8B",X"89",X"89",X"7F",
		X"74",X"74",X"74",X"75",X"76",X"77",X"78",X"78",X"7A",X"81",X"89",X"8D",X"8D",X"8C",X"8B",X"89",
		X"89",X"84",X"77",X"73",X"74",X"75",X"76",X"77",X"78",X"78",X"79",X"7E",X"86",X"8C",X"8D",X"8C",
		X"8C",X"8A",X"89",X"87",X"7C",X"74",X"74",X"75",X"76",X"76",X"77",X"78",X"78",X"7B",X"82",X"89",
		X"8D",X"8D",X"8C",X"8B",X"89",X"89",X"82",X"76",X"73",X"74",X"75",X"76",X"77",X"78",X"78",X"79",
		X"7E",X"86",X"8B",X"8D",X"8C",X"8B",X"8A",X"89",X"88",X"7C",X"74",X"74",X"75",X"75",X"76",X"77",
		X"78",X"78",X"7A",X"81",X"89",X"8C",X"8D",X"8C",X"8B",X"8A",X"8A",X"84",X"78",X"73",X"74",X"75",
		X"76",X"77",X"77",X"78",X"79",X"7C",X"84",X"8B",X"8D",X"8C",X"8B",X"8B",X"89",X"89",X"80",X"75",
		X"74",X"75",X"75",X"76",X"77",X"78",X"78",X"79",X"7E",X"86",X"8C",X"8D",X"8C",X"8B",X"8A",X"89",
		X"88",X"7C",X"74",X"74",X"75",X"75",X"76",X"77",X"78",X"78",X"7A",X"80",X"88",X"8C",X"8D",X"8C",
		X"8B",X"8A",X"8A",X"86",X"7A",X"74",X"74",X"75",X"76",X"76",X"77",X"78",X"79",X"7B",X"82",X"89",
		X"8C",X"8D",X"8B",X"8B",X"8A",X"89",X"84",X"78",X"74",X"74",X"75",X"76",X"77",X"77",X"78",X"79",
		X"7B",X"83",X"89",X"8C",X"8C",X"8B",X"8B",X"89",X"89",X"84",X"77",X"74",X"74",X"75",X"76",X"77",
		X"77",X"78",X"79",X"7C",X"83",X"8A",X"8C",X"8C",X"8B",X"8B",X"89",X"89",X"84",X"77",X"74",X"74",
		X"75",X"76",X"77",X"77",X"78",X"79",X"7B",X"82",X"89",X"8C",X"8C",X"8B",X"8B",X"89",X"89",X"84",
		X"77",X"74",X"74",X"75",X"76",X"77",X"78",X"78",X"79",X"7B",X"82",X"89",X"8C",X"8C",X"8B",X"8B",
		X"89",X"89",X"85",X"79",X"74",X"74",X"75",X"76",X"77",X"78",X"78",X"79",X"7B",X"81",X"88",X"8C",
		X"8C",X"8C",X"8B",X"8A",X"89",X"87",X"7B",X"74",X"74",X"75",X"76",X"77",X"77",X"78",X"79",X"7A",
		X"7F",X"86",X"8B",X"8C",X"8C",X"8B",X"8A",X"89",X"88",X"7E",X"75",X"74",X"75",X"76",X"76",X"77",
		X"78",X"79",X"79",X"7D",X"84",X"8A",X"8C",X"8C",X"8B",X"8A",X"89",X"89",X"82",X"76",X"74",X"74",
		X"76",X"76",X"77",X"78",X"79",X"79",X"7C",X"82",X"88",X"8C",X"8C",X"8B",X"8B",X"8A",X"89",X"85",
		X"79",X"74",X"75",X"75",X"76",X"77",X"78",X"78",X"79",X"7B",X"80",X"87",X"8B",X"8C",X"8C",X"8B",
		X"8A",X"89",X"87",X"7C",X"74",X"74",X"75",X"76",X"76",X"77",X"78",X"79",X"7A",X"7E",X"85",X"8A",
		X"8C",X"8C",X"8B",X"8A",X"89",X"89",X"7F",X"75",X"74",X"75",X"76",X"76",X"77",X"78",X"79",X"7A",
		X"7D",X"84",X"89",X"8C",X"8C",X"8B",X"8A",X"89",X"89",X"81",X"76",X"74",X"75",X"76",X"77",X"77",
		X"78",X"79",X"79",X"7D",X"83",X"89",X"8C",X"8C",X"8B",X"8A",X"89",X"89",X"81",X"76",X"74",X"75",
		X"76",X"77",X"77",X"78",X"79",X"7A",X"7D",X"83",X"89",X"8C",X"8C",X"8B",X"8A",X"89",X"89",X"80",
		X"75",X"74",X"75",X"76",X"77",X"78",X"78",X"79",X"7A",X"7E",X"84",X"89",X"8C",X"8C",X"8B",X"8A",
		X"89",X"88",X"7E",X"75",X"74",X"75",X"76",X"77",X"78",X"78",X"79",X"7B",X"7F",X"85",X"8A",X"8C",
		X"8C",X"8B",X"8A",X"89",X"86",X"7B",X"74",X"75",X"75",X"76",X"77",X"78",X"79",X"79",X"7B",X"80",
		X"87",X"8A",X"8C",X"8C",X"8B",X"89",X"89",X"84",X"78",X"74",X"75",X"75",X"76",X"77",X"78",X"79",
		X"7A",X"7C",X"82",X"88",X"8B",X"8C",X"8C",X"8B",X"89",X"89",X"80",X"76",X"74",X"75",X"76",X"77",
		X"78",X"79",X"79",X"7A",X"7E",X"85",X"8A",X"8C",X"8C",X"8B",X"8A",X"89",X"86",X"7A",X"74",X"75",
		X"75",X"77",X"77",X"78",X"79",X"7A",X"7C",X"82",X"87",X"8B",X"8C",X"8B",X"8B",X"89",X"89",X"80",
		X"75",X"75",X"75",X"76",X"77",X"78",X"78",X"79",X"7B",X"7F",X"85",X"89",X"8C",X"8C",X"8B",X"8A",
		X"8A",X"85",X"78",X"74",X"75",X"76",X"77",X"77",X"78",X"79",X"7A",X"7D",X"83",X"88",X"8B",X"8C",
		X"8B",X"8A",X"8A",X"87",X"7C",X"75",X"75",X"76",X"76",X"77",X"78",X"79",X"7A",X"7C",X"81",X"87",
		X"8A",X"8C",X"8C",X"8B",X"8A",X"89",X"7F",X"76",X"75",X"76",X"76",X"77",X"78",X"79",X"79",X"7B",
		X"80",X"86",X"89",X"8B",X"8C",X"8B",X"8A",X"89",X"81",X"77",X"75",X"76",X"76",X"77",X"78",X"79",
		X"79",X"7A",X"7F",X"85",X"89",X"8B",X"8B",X"8B",X"8A",X"8A",X"83",X"78",X"75",X"76",X"76",X"77",
		X"78",X"79",X"79",X"7A",X"7E",X"84",X"88",X"8B",X"8C",X"8B",X"8A",X"8A",X"84",X"78",X"75",X"76",
		X"76",X"77",X"78",X"79",X"79",X"7A",X"7E",X"84",X"88",X"8B",X"8C",X"8B",X"8A",X"89",X"83",X"78",
		X"75",X"76",X"76",X"77",X"78",X"79",X"79",X"7A",X"7E",X"84",X"88",X"8B",X"8C",X"8B",X"8A",X"8A",
		X"82",X"77",X"75",X"76",X"77",X"77",X"78",X"79",X"79",X"7B",X"7F",X"85",X"89",X"8B",X"8C",X"8B",
		X"8A",X"89",X"80",X"76",X"75",X"76",X"77",X"77",X"78",X"79",X"7A",X"7B",X"80",X"86",X"89",X"8B",
		X"8B",X"8B",X"8A",X"88",X"7D",X"76",X"75",X"76",X"77",X"78",X"78",X"79",X"7A",X"7C",X"82",X"86",
		X"8A",X"8B",X"8B",X"8A",X"8A",X"86",X"7A",X"75",X"76",X"76",X"77",X"78",X"79",X"79",X"7A",X"7E",
		X"83",X"88",X"8A",X"8B",X"8B",X"8A",X"8A",X"82",X"77",X"75",X"76",X"77",X"78",X"78",X"79",X"7A",
		X"7B",X"80",X"85",X"89",X"8B",X"8B",X"8B",X"8A",X"88",X"7D",X"76",X"76",X"76",X"77",X"78",X"79",
		X"79",X"7A",X"7D",X"82",X"87",X"8A",X"8B",X"8B",X"8A",X"8A",X"84",X"79",X"75",X"76",X"77",X"77",
		X"78",X"79",X"79",X"7B",X"7F",X"85",X"88",X"8A",X"8B",X"8B",X"8A",X"88",X"7D",X"76",X"76",X"76",
		X"77",X"78",X"79",X"79",X"7A",X"7D",X"82",X"87",X"8A",X"8B",X"8B",X"8A",X"8A",X"83",X"78",X"76",
		X"76",X"77",X"77",X"78",X"79",X"7A",X"7B",X"80",X"85",X"89",X"8A",X"8B",X"8A",X"8A",X"87",X"7B",
		X"76",X"76",X"77",X"77",X"78",X"79",X"79",X"7B",X"7E",X"84",X"88",X"8A",X"8B",X"8B",X"8A",X"89",
		X"7E",X"76",X"76",X"76",X"77",X"78",X"79",X"79",X"7A",X"7D",X"82",X"86",X"8A",X"8B",X"8B",X"8A",
		X"8A",X"81",X"77",X"76",X"76",X"77",X"78",X"79",X"79",X"7A",X"7C",X"81",X"86",X"89",X"8A",X"8B",
		X"8A",X"8A",X"84",X"78",X"76",X"76",X"77",X"78",X"79",X"79",X"7A",X"7B",X"80",X"85",X"88",X"8A",
		X"8B",X"8B",X"8A",X"85",X"7A",X"76",X"76",X"77",X"78",X"79",X"79",X"7A",X"7B",X"80",X"84",X"88",
		X"8A",X"8B",X"8B",X"8A",X"86",X"7B",X"76",X"76",X"77",X"78",X"79",X"7A",X"7A",X"7B",X"80",X"84",
		X"87",X"8A",X"8B",X"8B",X"8A",X"87",X"7B",X"76",X"76",X"77",X"78",X"79",X"79",X"7A",X"7B",X"7F",
		X"84",X"87",X"8A",X"8B",X"8A",X"8A",X"87",X"7B",X"76",X"77",X"77",X"78",X"79",X"79",X"7A",X"7B",
		X"80",X"84",X"87",X"8A",X"8B",X"8A",X"8B",X"86",X"7A",X"76",X"77",X"77",X"78",X"79",X"79",X"7A",
		X"7C",X"80",X"85",X"88",X"8A",X"8B",X"8A",X"8A",X"84",X"79",X"76",X"77",X"78",X"78",X"79",X"79",
		X"7A",X"7C",X"81",X"85",X"88",X"8A",X"8B",X"8A",X"8A",X"82",X"78",X"76",X"77",X"78",X"78",X"79",
		X"7A",X"7A",X"7D",X"82",X"86",X"88",X"8A",X"8B",X"8A",X"89",X"7F",X"77",X"77",X"77",X"78",X"78",
		X"79",X"7A",X"7B",X"7E",X"83",X"87",X"89",X"8A",X"8B",X"8A",X"87",X"7C",X"77",X"77",X"77",X"78",
		X"78",X"79",X"7A",X"7C",X"80",X"84",X"87",X"89",X"8A",X"8A",X"8A",X"84",X"7A",X"77",X"77",X"78",
		X"78",X"79",X"7A",X"7A",X"7D",X"81",X"85",X"88",X"8A",X"8A",X"8A",X"8A",X"81",X"78",X"77",X"77",
		X"78",X"78",X"79",X"7A",X"7A",X"7E",X"82",X"86",X"88",X"8A",X"8A",X"8A",X"88",X"7E",X"77",X"77",
		X"77",X"78",X"78",X"79",X"7A",X"7B",X"7F",X"83",X"87",X"89",X"8A",X"8A",X"8A",X"87",X"7C",X"77",
		X"77",X"78",X"78",X"79",X"79",X"7A",X"7B",X"80",X"84",X"87",X"89",X"8A",X"8A",X"8A",X"85",X"7A",
		X"77",X"77",X"78",X"79",X"79",X"7A",X"7A",X"7C",X"80",X"84",X"87",X"89",X"8A",X"8A",X"8A",X"85",
		X"7A",X"77",X"77",X"78",X"79",X"79",X"79",X"7A",X"7C",X"80",X"84",X"87",X"89",X"8A",X"8A",X"8A",
		X"84",X"7A",X"77",X"77",X"78",X"79",X"79",X"79",X"7A",X"7C",X"80",X"84",X"87",X"89",X"8A",X"8A",
		X"8A",X"85",X"7A",X"77",X"77",X"78",X"78",X"79",X"7A",X"7A",X"7C",X"80",X"84",X"86",X"88",X"8A",
		X"8A",X"8A",X"86",X"7B",X"77",X"77",X"78",X"78",X"79",X"7A",X"7A",X"7C",X"7F",X"83",X"86",X"88",
		X"89",X"8A",X"8A",X"87",X"7D",X"77",X"77",X"78",X"78",X"79",X"7A",X"7A",X"7B",X"7E",X"82",X"85",
		X"88",X"89",X"8A",X"8A",X"89",X"80",X"78",X"77",X"78",X"78",X"79",X"7A",X"7A",X"7B",X"7D",X"81",
		X"84",X"87",X"88",X"89",X"8A",X"89",X"83",X"79",X"77",X"78",X"78",X"79",X"7A",X"7A",X"7B",X"7C",
		X"80",X"83",X"86",X"88",X"89",X"89",X"89",X"86",X"7C",X"78",X"78",X"78",X"79",X"79",X"7A",X"7B",
		X"7B",X"7E",X"82",X"85",X"88",X"89",X"89",X"89",X"89",X"81",X"78",X"78",X"78",X"78",X"79",X"7A",
		X"7A",X"7B",X"7C",X"80",X"84",X"87",X"88",X"89",X"89",X"89",X"86",X"7C",X"77",X"78",X"78",X"79",
		X"79",X"7A",X"7A",X"7B",X"7E",X"82",X"85",X"88",X"89",X"89",X"89",X"89",X"81",X"78",X"78",X"78",
		X"79",X"79",X"7A",X"7A",X"7B",X"7C",X"80",X"83",X"86",X"88",X"89",X"89",X"89",X"87",X"7D",X"78",
		X"78",X"78",X"79",X"79",X"7A",X"7B",X"7B",X"7D",X"81",X"85",X"87",X"88",X"89",X"89",X"89",X"84",
		X"7A",X"78",X"78",X"78",X"79",X"7A",X"7A",X"7B",X"7B",X"7E",X"82",X"85",X"87",X"88",X"89",X"89",
		X"89",X"81",X"79",X"78",X"78",X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7F",X"83",X"86",X"87",X"88",
		X"89",X"89",X"88",X"7F",X"78",X"78",X"78",X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"80",X"84",X"86",
		X"87",X"88",X"89",X"89",X"87",X"7D",X"78",X"78",X"78",X"79",X"7A",X"7A",X"7B",X"7B",X"7D",X"80",
		X"84",X"86",X"87",X"88",X"88",X"89",X"86",X"7D",X"78",X"78",X"78",X"79",X"7A",X"7B",X"7B",X"7B",
		X"7D",X"80",X"84",X"86",X"87",X"88",X"88",X"89",X"86",X"7D",X"78",X"78",X"78",X"7A",X"7A",X"7B",
		X"7B",X"7B",X"7D",X"80",X"83",X"86",X"87",X"88",X"88",X"88",X"86",X"7D",X"78",X"78",X"79",X"7A",
		X"7A",X"7B",X"7B",X"7B",X"7D",X"80",X"83",X"86",X"87",X"88",X"88",X"88",X"87",X"7E",X"79",X"78",
		X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7D",X"80",X"83",X"85",X"87",X"87",X"88",X"88",X"87",X"80",
		X"79",X"78",X"79",X"79",X"7A",X"7B",X"7B",X"7C",X"7C",X"7F",X"83",X"85",X"86",X"87",X"88",X"88",
		X"88",X"81",X"79",X"78",X"79",X"79",X"7A",X"7B",X"7B",X"7C",X"7C",X"7F",X"82",X"85",X"86",X"87",
		X"88",X"88",X"88",X"81",X"79",X"78",X"78",X"79",X"7A",X"7B",X"7B",X"7C",X"7C",X"7F",X"82",X"85",
		X"86",X"87",X"88",X"88",X"88",X"82",X"79",X"78",X"78",X"79",X"7A",X"7B",X"7B",X"7C",X"7C",X"7F",
		X"82",X"85",X"86",X"87",X"88",X"88",X"88",X"81",X"79",X"78",X"78",X"79",X"7A",X"7B",X"7B",X"7C",
		X"7C",X"7F",X"83",X"85",X"86",X"87",X"88",X"88",X"87",X"80",X"79",X"78",X"79",X"7A",X"7A",X"7B",
		X"7B",X"7C",X"7D",X"80",X"83",X"85",X"86",X"87",X"88",X"88",X"87",X"7E",X"78",X"78",X"79",X"7A",
		X"7A",X"7B",X"7B",X"7C",X"7D",X"81",X"84",X"86",X"87",X"87",X"88",X"88",X"85",X"7C",X"78",X"79",
		X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7E",X"82",X"84",X"86",X"87",X"88",X"88",X"88",X"83",X"7A",
		X"78",X"79",X"79",X"7A",X"7B",X"7B",X"7B",X"7C",X"80",X"82",X"85",X"86",X"87",X"87",X"88",X"87",
		X"7F",X"79",X"79",X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7E",X"81",X"83",X"85",X"86",X"87",X"87",
		X"88",X"84",X"7B",X"79",X"79",X"79",X"7A",X"7B",X"7B",X"7B",X"7C",X"7F",X"82",X"84",X"86",X"87",
		X"87",X"88",X"87",X"7F",X"79",X"79",X"79",X"7A",X"7A",X"7B",X"7B",X"7C",X"7D",X"81",X"83",X"85",
		X"86",X"87",X"87",X"88",X"84",X"7B",X"79",X"79",X"7A",X"7A",X"7B",X"7B",X"7B",X"7C",X"80",X"83",
		X"84",X"86",X"87",X"87",X"87",X"86",X"7E",X"79",X"79",X"79",X"7A",X"7B",X"7B",X"7B",X"7C",X"7E",
		X"82",X"84",X"85",X"86",X"87",X"87",X"87",X"81",X"7A",X"79",X"79",X"7A",X"7B",X"7B",X"7B",X"7C",
		X"7D",X"81",X"83",X"85",X"86",X"87",X"87",X"88",X"83",X"7B",X"79",X"79",X"7A",X"7B",X"7B",X"7B",
		X"7C",X"7D",X"80",X"83",X"85",X"86",X"86",X"87",X"87",X"85",X"7C",X"79",X"79",X"7A",X"7B",X"7B",
		X"7B",X"7C",X"7D",X"7F",X"82",X"84",X"85",X"86",X"87",X"87",X"86",X"7E",X"79",X"7A",X"7A",X"7B",
		X"7B",X"7B",X"7C",X"7D",X"7F",X"82",X"84",X"85",X"86",X"87",X"87",X"86",X"7E",X"7A",X"7A",X"7A",
		X"7A",X"7B",X"7B",X"7B",X"7D",X"7F",X"82",X"84",X"85",X"86",X"86",X"87",X"86",X"7F",X"7A",X"7A",
		X"7A",X"7B",X"7B",X"7B",X"7C",X"7D",X"7F",X"82",X"84",X"85",X"86",X"86",X"87",X"86",X"7F",X"7A",
		X"7A",X"7A",X"7B",X"7B",X"7B",X"7C",X"7D",X"7F",X"82",X"84",X"85",X"86",X"86",X"87",X"86",X"7E",
		X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7C",X"7D",X"7F",X"82",X"84",X"85",X"86",X"86",X"87",X"85",
		X"7D",X"7A",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7D",X"80",X"82",X"84",X"85",X"86",X"86",X"87",
		X"84",X"7C",X"7A",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7E",X"80",X"82",X"84",X"85",X"86",X"86",
		X"87",X"82",X"7B",X"7A",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7E",X"81",X"83",X"85",X"85",X"86",
		X"86",X"86",X"80",X"7A",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7D",X"7F",X"81",X"84",X"85",X"86",
		X"86",X"87",X"85",X"7E",X"7A",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7D",X"80",X"82",X"84",X"85",
		X"86",X"86",X"86",X"83",X"7C",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7C",X"7E",X"81",X"83",X"84",
		X"85",X"86",X"86",X"86",X"80",X"7A",X"7A",X"7A",X"7B",X"7C",X"7C",X"7C",X"7D",X"7F",X"82",X"84",
		X"85",X"86",X"86",X"86",X"84",X"7D",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7C",X"7E",X"80",X"83",
		X"84",X"85",X"86",X"86",X"86",X"80",X"7B",X"7A",X"7A",X"7B",X"7C",X"7C",X"7C",X"7D",X"7F",X"81",
		X"83",X"85",X"85",X"86",X"86",X"83",X"7C",X"7A",X"7A",X"7B",X"7B",X"7C",X"7C",X"7D",X"7E",X"80",
		X"83",X"84",X"85",X"86",X"86",X"85",X"7F",X"7B",X"7A",X"7B",X"7B",X"7C",X"7C",X"7C",X"7E",X"80",
		X"82",X"83",X"85",X"85",X"86",X"86",X"81",X"7C",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7D",X"7F",
		X"81",X"83",X"84",X"85",X"85",X"86",X"83",X"7D",X"7B",X"7B",X"7B",X"7B",X"7C",X"7D",X"7D",X"7E",
		X"81",X"82",X"84",X"85",X"85",X"86",X"84",X"7F",X"7B",X"7B",X"7B",X"7B",X"7C",X"7D",X"7D",X"7E",
		X"80",X"82",X"83",X"85",X"85",X"85",X"85",X"80",X"7C",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",
		X"7F",X"81",X"83",X"84",X"85",X"85",X"86",X"82",X"7D",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",
		X"7F",X"80",X"82",X"84",X"85",X"85",X"86",X"84",X"7E",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7D",
		X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"85",X"80",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",
		X"7D",X"7F",X"81",X"83",X"84",X"85",X"85",X"86",X"83",X"7D",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",
		X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"85",X"80",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",
		X"7D",X"7D",X"7F",X"81",X"83",X"84",X"85",X"85",X"86",X"83",X"7D",X"7B",X"7B",X"7B",X"7C",X"7C",
		X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"85",X"81",X"7C",X"7B",X"7B",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7F",X"81",X"83",X"84",X"84",X"85",X"85",X"84",X"7F",X"7B",X"7B",X"7B",X"7C",
		X"7C",X"7C",X"7D",X"7D",X"7F",X"81",X"83",X"84",X"85",X"85",X"85",X"83",X"7E",X"7B",X"7B",X"7C",
		X"7C",X"7C",X"7C",X"7D",X"7E",X"7F",X"81",X"83",X"84",X"85",X"85",X"85",X"82",X"7D",X"7B",X"7B",
		X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"85",X"81",X"7C",X"7B",
		X"7B",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"85",X"81",X"7C",
		X"7B",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"85",X"80",
		X"7C",X"7B",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",X"85",
		X"80",X"7C",X"7B",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",X"85",
		X"85",X"81",X"7C",X"7B",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"85",
		X"85",X"85",X"82",X"7D",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"80",X"81",X"83",X"83",
		X"84",X"85",X"85",X"83",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7F",X"81",X"82",
		X"83",X"84",X"85",X"85",X"83",X"7F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7F",X"81",
		X"82",X"83",X"84",X"84",X"85",X"84",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",
		X"80",X"81",X"83",X"84",X"84",X"84",X"85",X"82",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",
		X"7D",X"7F",X"81",X"82",X"83",X"84",X"84",X"84",X"84",X"7F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",
		X"7D",X"7D",X"7E",X"80",X"82",X"83",X"84",X"84",X"84",X"84",X"82",X"7D",X"7C",X"7C",X"7C",X"7C",
		X"7D",X"7D",X"7D",X"7E",X"7F",X"81",X"82",X"83",X"84",X"84",X"84",X"84",X"80",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"80",X"81",X"83",X"83",X"84",X"84",X"84",X"82",X"7E",X"7C",
		X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7F",X"81",X"82",X"83",X"83",X"84",X"84",X"84",X"81",
		X"7D",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7F",X"81",X"82",X"83",X"84",X"84",X"84",
		X"84",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"80",X"81",X"82",X"83",X"84",
		X"84",X"84",X"83",X"7F",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"80",X"81",X"82",
		X"83",X"84",X"84",X"84",X"83",X"7E",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"80",
		X"81",X"82",X"83",X"84",X"84",X"84",X"82",X"7E",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",
		X"7F",X"80",X"81",X"82",X"83",X"84",X"84",X"84",X"83",X"7E",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7E",X"80",X"81",X"82",X"83",X"84",X"84",X"84",X"83",X"7F",X"7C",X"7C",X"7C",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7E",X"80",X"81",X"82",X"83",X"83",X"84",X"84",X"83",X"7F",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"80",X"81",X"82",X"83",X"83",X"84",X"84",X"83",X"80",
		X"7D",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7F",X"81",X"82",X"83",X"83",X"84",X"84",
		X"84",X"81",X"7D",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",
		X"83",X"84",X"84",X"82",X"7E",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"80",X"81",
		X"82",X"83",X"83",X"84",X"84",X"83",X"80",X"7D",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",
		X"7F",X"81",X"82",X"82",X"83",X"83",X"83",X"84",X"82",X"7E",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"83",X"83",X"84",X"83",X"7F",X"7C",X"7C",X"7C",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7E",X"7F",X"80",X"82",X"82",X"83",X"83",X"83",X"84",X"82",X"7E",X"7C",
		X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"80",X"81",X"82",X"82",X"83",X"83",X"83",X"83",
		X"80",X"7D",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"83",X"83",
		X"83",X"83",X"82",X"7F",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"82",
		X"82",X"83",X"83",X"83",X"83",X"82",X"7E",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",
		X"7F",X"81",X"82",X"82",X"83",X"83",X"83",X"83",X"81",X"7D",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",
		X"7E",X"7E",X"7E",X"80",X"81",X"82",X"82",X"83",X"83",X"83",X"83",X"81",X"7D",X"7C",X"7C",X"7D",
		X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"80",X"81",X"82",X"82",X"83",X"83",X"83",X"83",X"80",X"7D",
		X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",X"83",X"83",
		X"83",X"80",X"7D",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",
		X"83",X"83",X"83",X"83",X"81",X"7D",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"80",
		X"81",X"82",X"82",X"83",X"83",X"83",X"83",X"81",X"7D",X"7C",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",
		X"7E",X"7E",X"80",X"80",X"81",X"82",X"83",X"83",X"83",X"83",X"82",X"7E",X"7C",X"7D",X"7D",X"7D",
		X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"83",X"83",X"83",X"83",X"83",X"7F",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",X"83",X"83",
		X"83",X"80",X"7D",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"81",X"82",X"82",
		X"83",X"83",X"83",X"83",X"82",X"7E",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"80",X"81",X"82",X"82",X"83",X"83",X"83",X"82",X"80",X"7D",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",
		X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",X"82",X"83",X"83",X"83",X"82",X"7E",X"7C",X"7D",X"7D",
		X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",X"83",X"83",X"83",X"80",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",X"83",
		X"83",X"83",X"82",X"7F",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",
		X"81",X"82",X"82",X"83",X"83",X"83",X"82",X"7E",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"80",X"81",X"81",X"82",X"83",X"83",X"83",X"83",X"81",X"7E",X"7D",X"7D",X"7D",X"7D",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"83",X"83",X"83",X"83",X"81",X"7E",
		X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"82",X"83",
		X"83",X"82",X"81",X"7E",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",
		X"82",X"82",X"82",X"83",X"83",X"82",X"81",X"7E",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"80",X"81",X"82",X"82",X"82",X"83",X"83",X"83",X"81",X"7E",X"7D",X"7D",X"7D",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"81",X"7F",
		X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",
		X"82",X"83",X"82",X"7F",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",
		X"81",X"82",X"82",X"82",X"82",X"83",X"82",X"80",X"7E",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"83",X"81",X"7E",X"7D",X"7D",X"7D",
		X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"83",X"82",
		X"7F",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",
		X"82",X"82",X"82",X"82",X"81",X"7E",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"81",X"7F",X"7D",
		X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"82",X"82",X"82",X"82",
		X"82",X"82",X"81",X"7E",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"80",
		X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"7E",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"7E",X"7D",X"7D",
		X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"82",
		X"82",X"80",X"7E",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",
		X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"7E",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7F",X"7F",X"80",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"81",X"80",X"7E",X"7D",X"7D",X"7D",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"80",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"81",
		X"80",X"7E",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"81",X"81",X"81",
		X"82",X"82",X"82",X"82",X"81",X"80",X"7E",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"7F",X"80",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"81",X"80",X"7E",X"7D",X"7D",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"81",X"7F",
		X"7E",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"82",
		X"82",X"82",X"81",X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"80",
		X"80",X"81",X"81",X"81",X"81",X"82",X"81",X"81",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"7F",X"7F",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7F",X"7E",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",
		X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"7F",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",
		X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",
		X"81",X"81",X"81",X"81",X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"80",
		X"7F",X"7E",X"7E",X"7F",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"81",
		X"81",X"81",X"80",X"7F",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",X"7E",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"80",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"80",X"80",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"81",X"81",
		X"81",X"80",X"80",X"7F",X"7F",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"83",X"7F",X"AC",X"C9",X"C9",X"A2",X"57",X"4B",X"46",X"48",X"47",X"47",X"47",X"47",X"48",X"48",
		X"49",X"48",X"4A",X"45",X"3A",X"2E",X"23",X"1D",X"1E",X"1D",X"1E",X"1D",X"1D",X"1D",X"1D",X"1D",
		X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1B",X"1C",X"1B",X"1C",X"1B",X"1C",X"1B",X"1C",X"1B",X"1C",X"1B",
		X"1C",X"1B",X"1C",X"1B",X"1B",X"1B",X"1C",X"1B",X"1B",X"1B",X"1C",X"1C",X"1C",X"1C",X"1C",X"1D",
		X"1B",X"1D",X"1E",X"6D",X"C1",X"D2",X"D8",X"D6",X"D8",X"D7",X"D7",X"D5",X"D5",X"D4",X"D3",X"D3",
		X"D2",X"D2",X"D1",X"D0",X"CF",X"CF",X"CE",X"CD",X"CC",X"CC",X"CB",X"CB",X"CB",X"CA",X"C9",X"C9",
		X"C8",X"C8",X"C8",X"C7",X"C7",X"C6",X"C6",X"C5",X"C5",X"C4",X"C4",X"C3",X"C3",X"C2",X"C2",X"C2",
		X"C1",X"C1",X"C1",X"C0",X"C0",X"C0",X"BF",X"BF",X"BF",X"BE",X"BD",X"BD",X"BC",X"BC",X"BB",X"BB",
		X"BB",X"BB",X"BA",X"BA",X"BA",X"B9",X"B9",X"B8",X"B8",X"B8",X"B7",X"B7",X"B6",X"B6",X"B5",X"B5",
		X"B4",X"B4",X"B3",X"B3",X"B2",X"B2",X"B1",X"B1",X"B1",X"B0",X"B0",X"B0",X"AF",X"AF",X"AF",X"AF",
		X"AE",X"AE",X"AD",X"AD",X"AD",X"AD",X"AC",X"AC",X"AC",X"AC",X"AC",X"AB",X"AB",X"A6",X"9C",X"92",
		X"89",X"80",X"78",X"70",X"69",X"63",X"5D",X"57",X"52",X"4D",X"48",X"44",X"40",X"3D",X"39",X"36",
		X"32",X"2F",X"2B",X"2A",X"26",X"25",X"1F",X"38",X"87",X"AF",X"B6",X"B8",X"B8",X"B7",X"B6",X"B6",
		X"B5",X"B5",X"B4",X"B4",X"B3",X"B3",X"B3",X"B3",X"B2",X"B2",X"B1",X"B1",X"B0",X"B0",X"B0",X"AF",
		X"AF",X"AF",X"AE",X"AE",X"AE",X"AD",X"AD",X"AD",X"AC",X"AC",X"AC",X"AC",X"AC",X"AB",X"AB",X"AB",
		X"AB",X"AA",X"AA",X"AA",X"AA",X"A9",X"A9",X"A9",X"A8",X"A8",X"A8",X"A8",X"A7",X"A1",X"99",X"90",
		X"88",X"80",X"79",X"72",X"6C",X"66",X"61",X"5C",X"57",X"52",X"4E",X"4A",X"46",X"43",X"40",X"3E",
		X"3B",X"39",X"36",X"35",X"32",X"31",X"2C",X"4F",X"94",X"AD",X"B2",X"B2",X"B2",X"B2",X"B1",X"B1",
		X"B0",X"B0",X"B0",X"B0",X"AF",X"AF",X"AE",X"AE",X"AD",X"AD",X"AD",X"AD",X"AC",X"AC",X"AB",X"AB",
		X"AB",X"AB",X"AA",X"AA",X"A9",X"A9",X"A9",X"A9",X"A8",X"A8",X"A8",X"A8",X"A8",X"A7",X"A7",X"A7",
		X"A6",X"A6",X"A6",X"A5",X"A5",X"A5",X"A5",X"A4",X"A4",X"A4",X"A4",X"A4",X"A3",X"9D",X"95",X"8D",
		X"86",X"7F",X"79",X"73",X"6E",X"69",X"65",X"60",X"5C",X"58",X"55",X"51",X"4E",X"4C",X"49",X"46",
		X"43",X"41",X"3E",X"3D",X"3A",X"39",X"36",X"61",X"99",X"AA",X"AE",X"AE",X"AE",X"AD",X"AD",X"AD",
		X"AC",X"AC",X"AC",X"AC",X"AB",X"AB",X"AA",X"AA",X"AA",X"A9",X"A9",X"A9",X"A8",X"A8",X"A7",X"A7",
		X"A7",X"A7",X"A6",X"A6",X"A6",X"A6",X"A5",X"A5",X"A5",X"A5",X"A5",X"A4",X"A4",X"A4",X"A3",X"A3",
		X"A3",X"A3",X"A3",X"A3",X"A2",X"A2",X"A2",X"A2",X"A1",X"A1",X"A1",X"A1",X"A1",X"A1",X"A1",X"A0",
		X"A0",X"A0",X"9F",X"9F",X"9F",X"9F",X"9E",X"9E",X"9E",X"9E",X"9E",X"9D",X"9D",X"9D",X"9D",X"9D",
		X"9D",X"9D",X"9C",X"9C",X"9C",X"9B",X"9B",X"98",X"92",X"8B",X"85",X"7F",X"7A",X"75",X"70",X"6C",
		X"68",X"64",X"61",X"5D",X"5A",X"57",X"54",X"51",X"4F",X"4C",X"4A",X"47",X"45",X"43",X"41",X"3F",
		X"3E",X"3D",X"3C",X"3B",X"3A",X"39",X"37",X"36",X"35",X"34",X"33",X"32",X"30",X"2F",X"2E",X"2E",
		X"2D",X"2D",X"2D",X"2E",X"2E",X"2D",X"2D",X"2D",X"2D",X"2C",X"2C",X"2E",X"68",X"A7",X"B6",X"BB",
		X"BA",X"BB",X"B9",X"B9",X"B8",X"B8",X"B8",X"B8",X"B7",X"B7",X"B6",X"B6",X"B6",X"B5",X"B5",X"B4",
		X"B3",X"B2",X"B2",X"B2",X"B2",X"B1",X"B0",X"AA",X"A4",X"9F",X"9A",X"95",X"90",X"8B",X"87",X"83",
		X"7F",X"7B",X"77",X"74",X"71",X"6E",X"6B",X"68",X"66",X"64",X"62",X"60",X"5E",X"5C",X"5B",X"59",
		X"57",X"56",X"54",X"52",X"50",X"4F",X"4D",X"4C",X"4B",X"4A",X"49",X"49",X"48",X"48",X"47",X"46",
		X"46",X"46",X"45",X"45",X"44",X"43",X"42",X"42",X"40",X"41",X"3D",X"5C",X"A2",X"C0",X"C6",X"C7",
		X"C7",X"C6",X"C6",X"C5",X"C4",X"C4",X"C4",X"C3",X"C2",X"C2",X"C1",X"C1",X"C0",X"C0",X"BF",X"BF",
		X"BE",X"BE",X"BE",X"BE",X"BD",X"BD",X"BC",X"BC",X"BC",X"BB",X"BB",X"BA",X"BA",X"BA",X"B9",X"B9",
		X"B8",X"B8",X"B8",X"B7",X"B7",X"B7",X"B6",X"B6",X"B5",X"B5",X"B5",X"B4",X"B4",X"B4",X"B3",X"B3",
		X"B2",X"AE",X"A8",X"A3",X"9E",X"99",X"95",X"91",X"8D",X"89",X"86",X"82",X"7F",X"7C",X"79",X"76",
		X"73",X"71",X"6E",X"6C",X"6A",X"68",X"66",X"65",X"63",X"62",X"5F",X"7D",X"A7",X"B2",X"B5",X"B5",
		X"B5",X"B5",X"B4",X"B3",X"B3",X"B3",X"B2",X"B2",X"B1",X"B1",X"B0",X"B0",X"AF",X"AF",X"AE",X"AE",
		X"AD",X"AD",X"AC",X"AC",X"AB",X"AA",X"A7",X"A1",X"9C",X"97",X"93",X"8F",X"8B",X"87",X"83",X"7F",
		X"7C",X"79",X"76",X"72",X"6F",X"6C",X"69",X"66",X"63",X"61",X"5F",X"5D",X"5B",X"59",X"58",X"57",
		X"55",X"53",X"52",X"50",X"4F",X"4E",X"4C",X"4B",X"4A",X"48",X"47",X"46",X"45",X"43",X"43",X"41",
		X"42",X"42",X"42",X"40",X"40",X"3F",X"40",X"3E",X"3F",X"3B",X"4F",X"8A",X"A8",X"AE",X"AF",X"AE",
		X"AD",X"AC",X"AC",X"AB",X"AA",X"A9",X"A9",X"A8",X"A7",X"A6",X"A5",X"A5",X"A4",X"A3",X"A3",X"A2",
		X"A1",X"A0",X"A0",X"9F",X"9E",X"9E",X"9D",X"9D",X"9D",X"9D",X"9C",X"9C",X"9C",X"9C",X"9B",X"9B",
		X"9B",X"9B",X"9A",X"9A",X"99",X"99",X"99",X"99",X"98",X"98",X"98",X"98",X"98",X"97",X"97",X"97",
		X"93",X"8F",X"8A",X"86",X"82",X"7F",X"7B",X"78",X"75",X"72",X"6F",X"6C",X"6A",X"68",X"66",X"63",
		X"61",X"5F",X"5E",X"5C",X"5A",X"58",X"57",X"55",X"54",X"51",X"66",X"8C",X"98",X"9B",X"9B",X"9C",
		X"9B",X"9B",X"9B",X"9A",X"9A",X"9A",X"9A",X"99",X"99",X"99",X"98",X"98",X"97",X"97",X"97",X"96",
		X"96",X"96",X"95",X"95",X"95",X"95",X"95",X"95",X"94",X"94",X"94",X"94",X"93",X"93",X"93",X"93",
		X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8C",X"8B",X"8B",X"8B",X"8A",X"8A",
		X"8A",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"87",X"87",X"85",X"81",X"7D",X"7A",X"76",X"73",
		X"70",X"6D",X"6B",X"68",X"65",X"63",X"61",X"5F",X"5D",X"5B",X"59",X"57",X"55",X"54",X"53",X"51",
		X"51",X"4F",X"4F",X"4B",X"5B",X"7D",X"8B",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",
		X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8A",X"8A",X"8A",X"8A",X"88",
		X"84",X"81",X"7D",X"7A",X"77",X"74",X"71",X"6E",X"6C",X"69",X"67",X"64",X"62",X"60",X"5E",X"5C",
		X"5A",X"59",X"57",X"55",X"53",X"52",X"50",X"50",X"4C",X"59",X"7A",X"89",X"8C",X"8D",X"8D",X"8D",
		X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"8A",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"87",X"87",X"87",X"87",X"87",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"83",
		X"80",X"7D",X"7A",X"77",X"74",X"71",X"6E",X"6C",X"6A",X"67",X"65",X"63",X"61",X"5F",X"5D",X"5C",
		X"5A",X"58",X"57",X"55",X"54",X"52",X"51",X"50",X"4F",X"4E",X"4E",X"4D",X"4C",X"4B",X"4B",X"4A",
		X"49",X"48",X"47",X"47",X"46",X"46",X"45",X"45",X"44",X"44",X"44",X"44",X"44",X"45",X"45",X"45",
		X"45",X"46",X"43",X"57",X"82",X"94",X"98",X"99",X"99",X"99",X"98",X"98",X"97",X"97",X"97",X"97",
		X"97",X"97",X"96",X"96",X"96",X"96",X"95",X"95",X"95",X"95",X"94",X"95",X"94",X"94",X"94",X"94",
		X"94",X"93",X"93",X"93",X"93",X"93",X"92",X"92",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",
		X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",
		X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8A",X"8A",X"8A",
		X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"87",X"87",X"87",X"86",X"86",X"86",X"85",X"85",
		X"85",X"85",X"85",X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7D",X"7A",X"78",X"75",X"73",X"70",X"6E",
		X"6C",X"6A",X"68",X"66",X"64",X"62",X"61",X"5F",X"5E",X"5C",X"5B",X"5A",X"59",X"58",X"57",X"56",
		X"55",X"53",X"55",X"6C",X"7F",X"83",X"84",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"81",
		X"81",X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7D",X"7B",X"79",X"76",X"74",X"72",X"70",X"6E",X"6C",
		X"6A",X"68",X"67",X"65",X"63",X"62",X"60",X"5F",X"5E",X"5D",X"5C",X"5B",X"5A",X"59",X"58",X"57",
		X"56",X"55",X"55",X"55",X"54",X"53",X"53",X"52",X"51",X"51",X"50",X"50",X"4F",X"4F",X"4F",X"4F",
		X"4F",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4E",X"4D",X"4D",X"4D",X"66",X"85",X"8E",X"90",
		X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",
		X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",
		X"8D",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"89",X"89",X"86",X"84",X"81",X"7F",X"7D",X"7A",X"78",X"76",X"74",X"73",X"71",X"6F",X"6E",X"6C",
		X"6A",X"69",X"68",X"67",X"66",X"65",X"63",X"62",X"61",X"61",X"5E",X"62",X"77",X"85",X"88",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"85",X"83",X"81",X"7F",X"7D",X"7B",X"79",X"77",X"75",
		X"74",X"72",X"71",X"6F",X"6E",X"6D",X"6C",X"6A",X"6A",X"68",X"68",X"67",X"66",X"65",X"65",X"63",
		X"67",X"7C",X"89",X"8C",X"8D",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"8B",X"8A",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"85",X"83",X"81",X"7F",X"7D",X"7B",X"7A",X"78",X"76",X"75",
		X"73",X"72",X"71",X"70",X"6F",X"6D",X"6C",X"6B",X"6A",X"69",X"68",X"67",X"67",X"66",X"66",X"64",
		X"6F",X"82",X"89",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"89",X"89",X"89",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"86",X"87",
		X"86",X"86",X"85",X"85",X"84",X"84",X"83",X"81",X"7F",X"7D",X"7B",X"7A",X"79",X"77",X"76",X"75",
		X"73",X"72",X"70",X"6F",X"6E",X"6D",X"6C",X"6B",X"6A",X"69",X"69",X"68",X"67",X"67",X"66",X"65",
		X"64",X"64",X"63",X"63",X"62",X"62",X"61",X"61",X"61",X"60",X"60",X"60",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"5F",X"5E",X"5E",X"5E",X"5D",X"5E",X"5D",X"5E",X"5D",X"67",X"82",X"8E",X"91",X"91",X"91",
		X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"8C",X"8A",X"88",X"86",X"84",X"83",X"82",X"80",X"7F",X"7D",
		X"7C",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"72",X"71",X"71",X"70",X"70",X"6E",X"73",
		X"84",X"8E",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",X"8D",X"8C",X"8A",X"88",X"86",X"84",X"82",
		X"81",X"7F",X"7E",X"7D",X"7B",X"7A",X"78",X"77",X"76",X"75",X"73",X"72",X"71",X"70",X"6F",X"6E",
		X"6D",X"6C",X"6C",X"6B",X"6A",X"6A",X"69",X"69",X"68",X"68",X"67",X"67",X"67",X"66",X"66",X"65",
		X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"65",X"64",X"64",X"63",X"64",X"64",X"64",X"64",X"74",
		X"8B",X"92",X"94",X"94",X"94",X"94",X"94",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"92",X"92",
		X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",
		X"8E",X"8E",X"8E",X"8D",X"8D",X"8B",X"89",X"88",X"86",X"84",X"83",X"81",X"80",X"7F",X"7E",X"7C",
		X"7B",X"7A",X"79",X"78",X"77",X"76",X"75",X"74",X"73",X"72",X"72",X"71",X"71",X"70",X"70",X"6F",
		X"6F",X"6E",X"6E",X"6D",X"6D",X"6D",X"6C",X"6C",X"6B",X"6B",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",
		X"6A",X"6A",X"6A",X"6A",X"69",X"6A",X"69",X"6A",X"69",X"76",X"8B",X"93",X"95",X"95",X"95",X"95",
		X"95",X"94",X"94",X"94",X"94",X"94",X"94",X"94",X"93",X"93",X"93",X"93",X"92",X"92",X"92",X"91",
		X"91",X"91",X"91",X"91",X"90",X"8E",X"8C",X"8B",X"89",X"88",X"86",X"85",X"84",X"82",X"81",X"80",
		X"7F",X"7D",X"7C",X"7B",X"7B",X"7A",X"79",X"78",X"78",X"77",X"76",X"76",X"75",X"74",X"7B",X"89",
		X"8F",X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",
		X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",
		X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8A",X"8A",X"8A",
		X"8A",X"8A",X"89",X"89",X"88",X"87",X"85",X"83",X"82",X"80",X"7F",X"7E",X"7D",X"7B",X"7A",X"79",
		X"78",X"77",X"76",X"75",X"74",X"74",X"73",X"72",X"71",X"70",X"6F",X"6F",X"6E",X"6D",X"6D",X"6D",
		X"6D",X"6C",X"6C",X"6B",X"6B",X"6A",X"6A",X"6A",X"6A",X"69",X"69",X"69",X"68",X"68",X"68",X"68",
		X"68",X"68",X"68",X"68",X"68",X"68",X"68",X"67",X"67",X"67",X"68",X"68",X"68",X"68",X"67",X"67",
		X"67",X"67",X"67",X"67",X"68",X"68",X"68",X"68",X"68",X"68",X"68",X"68",X"68",X"69",X"69",X"69",
		X"69",X"69",X"69",X"69",X"69",X"69",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",
		X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6E",X"6D",X"71",X"87",X"98",
		X"9C",X"9D",X"9D",X"9D",X"9D",X"9C",X"9C",X"9C",X"9C",X"9C",X"9B",X"9B",X"9B",X"9A",X"9A",X"9A",
		X"9A",X"99",X"99",X"99",X"99",X"98",X"98",X"98",X"97",X"96",X"94",X"93",X"92",X"90",X"8F",X"8D",
		X"8C",X"8B",X"89",X"88",X"86",X"85",X"84",X"83",X"82",X"82",X"81",X"80",X"7F",X"7E",X"7E",X"7E",
		X"7D",X"7C",X"80",X"8D",X"94",X"95",X"95",X"95",X"95",X"94",X"94",X"94",X"94",X"94",X"94",X"94",
		X"93",X"93",X"93",X"93",X"93",X"92",X"92",X"92",X"92",X"92",X"91",X"91",X"91",X"90",X"8F",X"8E",
		X"8C",X"8B",X"8A",X"88",X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"80",X"7F",X"7E",X"7D",X"7C",
		X"7C",X"7B",X"7A",X"7A",X"79",X"79",X"78",X"77",X"77",X"77",X"76",X"76",X"75",X"75",X"75",X"74",
		X"74",X"74",X"73",X"73",X"73",X"72",X"72",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"70",
		X"71",X"70",X"7A",X"8C",X"92",X"93",X"94",X"94",X"93",X"93",X"93",X"93",X"93",X"92",X"92",X"92",
		X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",
		X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",
		X"8B",X"8B",X"8B",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",
		X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"87",X"86",X"86",X"86",X"86",X"86",X"86",
		X"86",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"84",X"84",X"84",X"82",X"81",X"80",
		X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"78",X"77",X"77",X"76",X"75",X"74",X"74",X"73",X"73",
		X"72",X"72",X"71",X"71",X"71",X"70",X"72",X"7C",X"83",X"85",X"85",X"85",X"85",X"85",X"85",X"85",
		X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"84",X"84",X"84",X"84",X"84",X"84",
		X"84",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
		X"83",X"83",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"82",X"82",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",X"7E",X"7D",X"7C",X"7B",X"7A",X"79",X"78",X"78",
		X"77",X"76",X"75",X"74",X"74",X"73",X"72",X"72",X"71",X"70",X"70",X"6F",X"6F",X"6E",X"6E",X"6D",
		X"6D",X"6D",X"6C",X"6C",X"6C",X"6B",X"6B",X"6B",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",
		X"6A",X"69",X"69",X"69",X"69",X"6A",X"6A",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",
		X"69",X"69",X"69",X"69",X"69",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6A",X"6A",
		X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6C",
		X"6D",X"6C",X"6D",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6F",X"6F",X"6F",X"6F",X"70",X"6F",
		X"72",X"83",X"8F",X"91",X"92",X"92",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"91",X"91",
		X"91",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"8D",X"8C",X"8B",X"8A",
		X"89",X"88",X"87",X"86",X"85",X"84",X"83",X"82",X"82",X"81",X"80",X"80",X"7F",X"7F",X"7E",X"7E",
		X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"85",X"8C",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",
		X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"8B",X"8A",X"89",X"88",X"87",X"86",X"85",X"84",X"83",X"83",X"82",X"81",X"80",X"80",X"7F",X"7E",
		X"7D",X"7D",X"7C",X"7C",X"7B",X"7B",X"7A",X"7A",X"79",X"79",X"79",X"78",X"78",X"78",X"77",X"77",
		X"77",X"77",X"76",X"76",X"76",X"76",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"74",X"74",X"74",
		X"74",X"74",X"74",X"74",X"73",X"78",X"85",X"8B",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",
		X"8D",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"8A",X"89",X"88",X"87",X"86",X"85",X"84",X"83",X"82",X"81",X"80",X"80",X"7F",X"7E",X"7E",X"7D",
		X"7D",X"7C",X"7C",X"7B",X"7A",X"7A",X"79",X"79",X"78",X"78",X"78",X"78",X"77",X"77",X"77",X"76",
		X"76",X"76",X"75",X"75",X"75",X"75",X"74",X"74",X"74",X"74",X"73",X"73",X"73",X"73",X"73",X"73",
		X"72",X"72",X"72",X"72",X"72",X"72",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"70",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"72",
		X"72",X"72",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"76",
		X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"78",X"78",X"78",X"78",X"79",X"79",X"79",X"79",X"79",X"78",X"78",X"78",X"7B",X"8A",
		X"95",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"99",X"99",X"99",X"98",X"98",X"97",X"97",X"97",
		X"97",X"96",X"96",X"96",X"96",X"96",X"95",X"95",X"95",X"95",X"95",X"94",X"94",X"94",X"94",X"94",
		X"93",X"93",X"93",X"93",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",
		X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8A",
		X"8A",X"89",X"88",X"87",X"86",X"86",X"85",X"84",X"83",X"82",X"82",X"81",X"81",X"80",X"7F",X"7F",
		X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"82",X"89",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",
		X"89",X"88",X"88",X"88",X"87",X"87",X"86",X"85",X"84",X"83",X"83",X"82",X"81",X"80",X"80",X"7F",
		X"7F",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7B",X"7B",X"7B",X"7A",X"7A",X"79",X"79",X"78",X"78",
		X"78",X"78",X"78",X"78",X"77",X"77",X"77",X"77",X"76",X"76",X"76",X"76",X"76",X"75",X"75",X"75",
		X"74",X"74",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",
		X"74",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"74",
		X"74",X"74",X"75",X"7E",X"89",X"8C",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",
		X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8A",X"8A",X"89",
		X"88",X"87",X"87",X"86",X"85",X"85",X"84",X"83",X"83",X"82",X"81",X"81",X"80",X"80",X"7F",X"7E",
		X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"80",X"87",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"87",
		X"87",X"87",X"87",X"86",X"85",X"85",X"84",X"83",X"83",X"82",X"81",X"81",X"80",X"7F",X"7E",X"7E",
		X"7D",X"7D",X"7C",X"7C",X"7B",X"7B",X"7A",X"7A",X"7A",X"7A",X"79",X"79",X"78",X"7B",X"82",X"85",
		X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"84",
		X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"83",X"83",X"82",X"81",X"81",X"80",X"7F",X"7E",X"7E",
		X"7D",X"7C",X"7C",X"7B",X"7B",X"7A",X"79",X"78",X"77",X"77",X"76",X"76",X"76",X"76",X"76",X"75",
		X"75",X"75",X"78",X"7F",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"7F",
		X"7F",X"7E",X"7D",X"7C",X"7C",X"7B",X"7B",X"7A",X"7A",X"79",X"79",X"79",X"78",X"78",X"77",X"77",
		X"76",X"76",X"76",X"75",X"75",X"75",X"75",X"74",X"74",X"74",X"74",X"74",X"73",X"73",X"73",X"73",
		X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"72",X"72",X"72",X"72",X"71",X"71",X"71",X"71",X"71",
		X"71",X"72",X"79",X"81",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"83",
		X"83",X"83",X"84",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"81",
		X"80",X"7F",X"7F",X"7E",X"7E",X"7D",X"7D",X"7D",X"7C",X"7C",X"7B",X"7B",X"7B",X"7A",X"7D",X"89",
		X"97",X"A4",X"AC",X"AF",X"B0",X"B0",X"AF",X"A9",X"9A",X"8B",X"83",X"81",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7E",X"7E",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7D",X"84",X"90",X"9B",X"A3",X"A7",X"A8",X"A8",X"A8",X"A7",
		X"A6",X"A6",X"A5",X"A5",X"A4",X"A4",X"A3",X"A3",X"A3",X"A2",X"A2",X"A2",X"A1",X"A1",X"A0",X"A0",
		X"9F",X"9F",X"9E",X"9D",X"9D",X"9C",X"9C",X"9C",X"9B",X"9B",X"9A",X"9A",X"9A",X"9A",X"99",X"99",
		X"98",X"98",X"98",X"97",X"96",X"96",X"95",X"95",X"95",X"94",X"94",X"92",X"86",X"75",X"6A",X"66",
		X"65",X"65",X"66",X"66",X"66",X"66",X"66",X"66",X"67",X"67",X"67",X"67",X"67",X"67",X"67",X"68",
		X"68",X"68",X"68",X"68",X"68",X"68",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"69",X"6A",
		X"6A",X"6A",X"6A",X"6A",X"6B",X"6A",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",X"6B",
		X"6B",X"70",X"7B",X"84",X"8D",X"93",X"96",X"98",X"98",X"98",X"97",X"97",X"97",X"96",X"96",X"95",
		X"95",X"95",X"94",X"94",X"94",X"93",X"93",X"93",X"93",X"92",X"92",X"92",X"92",X"92",X"92",X"91",
		X"91",X"90",X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",
		X"8D",X"8D",X"8D",X"8C",X"8C",X"8A",X"7C",X"6A",X"62",X"5F",X"5F",X"5E",X"5F",X"5F",X"60",X"60",
		X"60",X"60",X"60",X"61",X"61",X"61",X"61",X"62",X"62",X"62",X"62",X"63",X"63",X"63",X"63",X"63",
		X"63",X"64",X"64",X"64",X"64",X"65",X"65",X"65",X"65",X"65",X"66",X"66",X"66",X"66",X"66",X"67",
		X"67",X"67",X"67",X"67",X"68",X"68",X"68",X"69",X"69",X"69",X"69",X"6E",X"77",X"7F",X"87",X"8D",
		X"91",X"94",X"95",X"95",X"94",X"94",X"94",X"94",X"94",X"93",X"93",X"93",X"93",X"92",X"92",X"92",
		X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",
		X"8E",X"8E",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"8B",X"8B",X"8A",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"87",
		X"87",X"87",X"88",X"87",X"87",X"87",X"87",X"87",X"86",X"86",X"86",X"85",X"85",X"85",X"84",X"84",
		X"84",X"84",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"81",X"81",
		X"81",X"81",X"81",X"80",X"80",X"77",X"65",X"59",X"56",X"55",X"55",X"55",X"56",X"56",X"57",X"57",
		X"57",X"57",X"58",X"58",X"59",X"59",X"5A",X"5A",X"5B",X"5B",X"5C",X"5C",X"5D",X"5D",X"5D",X"5F",
		X"65",X"6C",X"73",X"79",X"7F",X"83",X"86",X"88",X"88",X"89",X"89",X"89",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"87",X"87",X"87",X"87",X"87",X"86",X"86",X"86",X"86",X"86",X"86",X"86",
		X"86",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"84",X"84",X"84",X"84",X"83",X"84",
		X"83",X"83",X"83",X"83",X"7F",X"6F",X"5F",X"5A",X"58",X"59",X"59",X"59",X"59",X"5A",X"5A",X"5A",
		X"5A",X"5B",X"5B",X"5C",X"5C",X"5C",X"5C",X"5D",X"5D",X"5E",X"5E",X"5E",X"5E",X"5F",X"5F",X"5F",
		X"5F",X"60",X"60",X"60",X"61",X"61",X"61",X"62",X"62",X"62",X"63",X"63",X"63",X"63",X"64",X"64",
		X"64",X"64",X"65",X"65",X"65",X"65",X"66",X"66",X"66",X"66",X"67",X"67",X"67",X"68",X"68",X"68",
		X"68",X"69",X"69",X"69",X"69",X"69",X"69",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",
		X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6E",X"6F",
		X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"71",
		X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"72",X"73",X"73",X"74",X"74",X"74",X"74",X"74",X"74",
		X"74",X"74",X"74",X"75",X"75",X"75",X"75",X"75",X"76",X"77",X"7C",X"81",X"86",X"8A",X"8E",X"92",
		X"95",X"98",X"9A",X"9C",X"9D",X"9E",X"9E",X"9D",X"9D",X"9D",X"9D",X"9C",X"9C",X"9C",X"9B",X"9B",
		X"9B",X"9A",X"9A",X"9A",X"9A",X"9A",X"9A",X"99",X"99",X"99",X"99",X"98",X"98",X"98",X"98",X"98",
		X"97",X"97",X"97",X"96",X"96",X"96",X"95",X"95",X"95",X"95",X"94",X"94",X"94",X"94",X"8F",X"7C",
		X"6F",X"6B",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",
		X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"71",X"75",X"7A",X"7F",X"83",X"87",X"8A",
		X"8D",X"90",X"93",X"95",X"96",X"97",X"97",X"98",X"98",X"97",X"97",X"96",X"96",X"96",X"96",X"95",
		X"95",X"94",X"95",X"91",X"80",X"71",X"6D",X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",
		X"6C",X"6D",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6F",X"6F",X"6F",X"6F",X"6F",X"71",X"75",
		X"79",X"7E",X"81",X"85",X"88",X"8B",X"8E",X"90",X"93",X"94",X"95",X"96",X"97",X"97",X"97",X"97",
		X"97",X"97",X"96",X"96",X"95",X"95",X"94",X"94",X"91",X"80",X"71",X"6C",X"6B",X"6B",X"6B",X"6C",
		X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"71",X"71",
		X"71",X"71",X"72",X"73",X"77",X"7B",X"7F",X"83",X"86",X"89",X"8C",X"8F",X"91",X"94",X"95",X"97",
		X"98",X"98",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"98",X"98",X"97",
		X"97",X"97",X"96",X"96",X"96",X"96",X"95",X"95",X"95",X"95",X"95",X"94",X"94",X"94",X"94",X"93",
		X"93",X"93",X"93",X"92",X"92",X"92",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"91",X"90",
		X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",
		X"8D",X"8D",X"8B",X"7C",X"6C",X"66",X"65",X"65",X"65",X"66",X"66",X"67",X"67",X"67",X"67",X"67",
		X"68",X"68",X"68",X"69",X"69",X"69",X"69",X"6A",X"6A",X"6A",X"6B",X"6B",X"6C",X"6D",X"70",X"74",
		X"77",X"7A",X"7E",X"81",X"83",X"86",X"88",X"8A",X"8C",X"8E",X"8F",X"90",X"91",X"92",X"93",X"93",
		X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"92",X"92",X"92",X"91",
		X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",
		X"8C",X"8D",X"87",X"75",X"69",X"66",X"66",X"66",X"66",X"67",X"67",X"67",X"67",X"67",X"67",X"67",
		X"68",X"68",X"68",X"69",X"69",X"6A",X"6A",X"6A",X"6A",X"6B",X"6B",X"6B",X"6C",X"6D",X"71",X"74",
		X"77",X"7A",X"7D",X"7F",X"82",X"84",X"86",X"88",X"8A",X"8C",X"8D",X"8E",X"8F",X"90",X"91",X"91",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",X"91",X"91",X"91",
		X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8E",X"8E",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",
		X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8C",X"88",X"78",X"6A",X"67",
		X"66",X"66",X"66",X"67",X"67",X"67",X"67",X"68",X"68",X"68",X"68",X"68",X"69",X"69",X"69",X"6A",
		X"6B",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6D",X"70",X"73",X"76",X"79",X"7B",X"7D",X"7F",X"81",
		X"83",X"85",X"87",X"88",X"8A",X"8B",X"8C",X"8D",X"8D",X"8E",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"90",X"8E",X"80",X"71",X"6C",X"6B",X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6D",X"6C",X"6D",X"6C",
		X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",X"6F",X"6F",X"70",X"70",X"71",X"71",
		X"71",X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",X"78",X"78",
		X"78",X"78",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7D",X"80",X"82",X"84",
		X"86",X"88",X"89",X"8B",X"8C",X"8E",X"8F",X"90",X"91",X"92",X"93",X"94",X"94",X"95",X"96",X"96",
		X"97",X"97",X"98",X"98",X"98",X"98",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"98",
		X"98",X"98",X"98",X"98",X"98",X"97",X"97",X"97",X"97",X"96",X"96",X"96",X"96",X"95",X"95",X"95",
		X"95",X"95",X"94",X"94",X"94",X"94",X"94",X"94",X"93",X"93",X"93",X"93",X"93",X"92",X"92",X"92",
		X"92",X"91",X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",
		X"8B",X"8B",X"8B",X"8B",X"8C",X"86",X"76",X"6C",X"69",X"69",X"69",X"69",X"6A",X"6A",X"6A",X"6B",
		X"6B",X"6B",X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",X"6E",
		X"6F",X"6F",X"6F",X"6F",X"6F",X"6F",X"70",X"70",X"70",X"70",X"70",X"70",X"71",X"71",X"71",X"71",
		X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"72",X"73",X"73",X"73",X"74",X"77",X"79",X"7B",X"7D",
		X"7E",X"80",X"81",X"83",X"84",X"85",X"87",X"88",X"88",X"89",X"8A",X"8B",X"8C",X"8C",X"8D",X"8D",
		X"8E",X"8E",X"8F",X"8F",X"8F",X"90",X"90",X"90",X"91",X"91",X"91",X"91",X"91",X"91",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8E",X"8D",
		X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"86",X"77",X"6E",X"6C",X"6B",X"6B",
		X"6B",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6C",X"6D",X"6D",X"6D",X"6D",X"6D",X"6E",X"6E",X"6E",
		X"6E",X"6F",X"6F",X"6F",X"6F",X"70",X"72",X"74",X"75",X"77",X"79",X"7A",X"7B",X"7C",X"7D",X"7E",
		X"80",X"81",X"82",X"83",X"84",X"84",X"85",X"86",X"86",X"87",X"88",X"88",X"88",X"89",X"89",X"7F",
		X"74",X"71",X"70",X"70",X"70",X"71",X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",
		X"72",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"75",
		X"75",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",X"78",X"78",
		X"78",X"78",X"78",X"78",X"79",X"7B",X"7C",X"7E",X"80",X"81",X"82",X"83",X"84",X"86",X"86",X"87",
		X"88",X"89",X"8A",X"8A",X"8B",X"8B",X"8C",X"8C",X"8C",X"8D",X"8D",X"8D",X"8D",X"8E",X"8C",X"82",
		X"7A",X"78",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",X"78",
		X"78",X"78",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"81",X"82",X"82",X"83",X"84",X"85",X"86",X"87",X"88",X"89",X"8A",X"8A",X"8B",X"8C",X"8D",X"8E",
		X"8E",X"8E",X"8F",X"8F",X"8F",X"90",X"90",X"90",X"90",X"91",X"91",X"91",X"91",X"91",X"92",X"92",
		X"92",X"92",X"92",X"92",X"92",X"92",X"93",X"93",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",
		X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"91",X"91",X"91",X"91",X"91",
		X"91",X"91",X"91",X"91",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"8F",X"8F",X"8F",X"8F",X"8E",X"8E",X"8E",X"8E",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8C",
		X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",X"8B",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",
		X"8A",X"8A",X"8A",X"89",X"89",X"89",X"89",X"89",X"89",X"89",X"88",X"88",X"88",X"88",X"88",X"87",
		X"87",X"87",X"87",X"7E",X"74",X"71",X"70",X"70",X"6F",X"70",X"70",X"70",X"70",X"70",X"70",X"70",
		X"70",X"71",X"71",X"71",X"71",X"71",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",
		X"72",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"74",X"74",
		X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"73",X"73",X"74",X"74",X"74",X"74",X"75",X"75",
		X"75",X"75",X"75",X"75",X"75",X"75",X"75",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",
		X"76",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"78",X"78",X"78",X"78",X"78",X"78",
		X"78",X"78",X"78",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"7A",X"7C",
		X"7D",X"7E",X"7F",X"80",X"80",X"81",X"82",X"83",X"83",X"84",X"84",X"85",X"85",X"86",X"86",X"86",
		X"87",X"87",X"87",X"87",X"87",X"87",X"88",X"86",X"7F",X"7A",X"79",X"79",X"79",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"83",X"83",X"84",X"85",X"86",X"86",X"87",
		X"87",X"88",X"88",X"88",X"89",X"89",X"89",X"8A",X"8A",X"8A",X"8A",X"8B",X"8B",X"8B",X"8B",X"8B",
		X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",
		X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8B",X"8B",X"8B",X"8B",
		X"8B",X"8B",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"89",X"89",X"89",
		X"89",X"89",X"89",X"88",X"88",X"88",X"86",X"80",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7D",X"7D",X"7E",
		X"7F",X"80",X"80",X"81",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"83",X"83",X"83",X"83",X"84",
		X"84",X"84",X"84",X"84",X"84",X"84",X"81",X"7D",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7F",X"7F",X"80",
		X"80",X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"83",X"83",X"83",X"83",X"83",X"84",X"84",X"84",
		X"84",X"84",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"84",X"84",X"85",X"85",X"85",
		X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"85",X"84",X"84",X"84",X"84",X"84",
		X"81",X"7C",X"7B",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",
		X"83",X"83",X"83",X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"84",X"85",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"83",
		X"7E",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7E",X"7E",X"7F",
		X"7F",X"80",X"80",X"80",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"83",X"83",X"83",X"83",X"83",
		X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"84",X"83",X"84",X"83",
		X"83",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"82",X"7E",X"7B",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"79",X"79",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"7D",X"7C",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",
		X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"82",X"81",X"7E",X"7C",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7A",X"7A",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",X"7B",
		X"7B",X"7B",X"7B",X"7B",X"7B",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"81",X"81",X"81",
		X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"83",X"83",X"83",X"82",X"83",
		X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"81",X"7F",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7D",X"7D",X"7D",X"7D",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"81",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",
		X"7F",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"83",X"83",X"83",X"83",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"81",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"82",X"82",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"82",X"82",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"80",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"81",X"80",X"80",X"80",X"81",X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"80",X"7F",
		X"80",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",
		X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",
		X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",
		X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"7F",
		X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",
		X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"80",
		X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"7F",
		X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",
		X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",
		X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",
		X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"7F",X"80",
		X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",
		X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",
		X"7F",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",
		X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",
		X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",
		X"80",X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",
		X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",
		X"7F",X"80",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"80",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",
		X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"7F",
		X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",
		X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"80",
		X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",
		X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",
		X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",
		X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",
		X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"7F",
		X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",
		X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"80",
		X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",
		X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",
		X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",
		X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",
		X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",
		X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",
		X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",
		X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",
		X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",
		X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",
		X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"80",
		X"7F",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",
		X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"7F",
		X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",
		X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"7F",
		X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",
		X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",
		X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",
		X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",
		X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",
		X"80",X"7F",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",
		X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",
		X"7C",X"BA",X"A6",X"70",X"88",X"C5",X"DA",X"B6",X"7F",X"76",X"B7",X"DA",X"C8",X"8C",X"6E",X"9E",
		X"D7",X"D2",X"9E",X"6C",X"87",X"C8",X"D9",X"AF",X"73",X"74",X"B4",X"DC",X"C2",X"83",X"69",X"9E",
		X"D6",X"D0",X"95",X"67",X"85",X"C7",X"D9",X"A8",X"6C",X"72",X"B3",X"D9",X"BA",X"79",X"66",X"9C",
		X"D4",X"CB",X"8D",X"62",X"86",X"C6",X"D5",X"A1",X"66",X"70",X"B1",X"D6",X"B5",X"72",X"62",X"9A",
		X"D0",X"C6",X"85",X"5E",X"84",X"C4",X"D1",X"9C",X"62",X"6E",X"AF",X"D2",X"B0",X"6D",X"5F",X"97",
		X"CC",X"C1",X"81",X"59",X"7E",X"BF",X"CD",X"98",X"5E",X"6A",X"AB",X"CF",X"AD",X"6A",X"5A",X"92",
		X"C8",X"BE",X"7E",X"55",X"7A",X"BA",X"C9",X"95",X"5A",X"65",X"A6",X"CC",X"AC",X"68",X"57",X"8E",
		X"C5",X"BC",X"7C",X"52",X"75",X"B6",X"C6",X"94",X"58",X"60",X"A0",X"C8",X"AA",X"68",X"53",X"88",
		X"C1",X"BC",X"7E",X"50",X"6E",X"B0",X"C5",X"96",X"57",X"5A",X"99",X"C4",X"AC",X"69",X"4E",X"7F",
		X"BB",X"BC",X"81",X"4E",X"67",X"A9",X"C3",X"99",X"58",X"53",X"90",X"C1",X"AE",X"6C",X"4A",X"76",
		X"B4",X"BD",X"86",X"4E",X"5E",X"A0",X"C2",X"A0",X"5D",X"4D",X"84",X"BB",X"B2",X"72",X"48",X"6A",
		X"AB",X"BD",X"8C",X"4F",X"55",X"95",X"BF",X"A5",X"63",X"49",X"7B",X"B6",X"B6",X"7B",X"48",X"61",
		X"A2",X"BE",X"95",X"55",X"4D",X"88",X"BB",X"AC",X"6B",X"45",X"6C",X"AB",X"BA",X"87",X"4B",X"53",
		X"93",X"BC",X"A0",X"5D",X"45",X"77",X"B2",X"B3",X"77",X"45",X"5C",X"9E",X"BB",X"93",X"52",X"49",
		X"83",X"B6",X"A9",X"69",X"42",X"67",X"A7",X"B7",X"85",X"49",X"4F",X"8F",X"B9",X"9F",X"5D",X"43",
		X"74",X"AF",X"B2",X"77",X"43",X"58",X"9A",X"B9",X"93",X"51",X"46",X"7F",X"B4",X"AA",X"6B",X"41",
		X"63",X"A3",X"B7",X"88",X"4A",X"4B",X"89",X"B7",X"A2",X"60",X"40",X"6B",X"A9",X"B3",X"7D",X"44",
		X"51",X"91",X"B7",X"99",X"57",X"41",X"74",X"AE",X"AE",X"72",X"40",X"57",X"98",X"B6",X"8F",X"4E",
		X"43",X"7C",X"B1",X"A8",X"68",X"3E",X"5F",X"A0",X"B5",X"87",X"48",X"47",X"84",X"B3",X"A1",X"60",
		X"3D",X"65",X"A4",X"B2",X"7F",X"44",X"4B",X"8B",X"B5",X"9C",X"5A",X"3E",X"6C",X"A9",X"B0",X"78",
		X"41",X"50",X"90",X"B5",X"96",X"54",X"3E",X"71",X"AC",X"AD",X"72",X"3F",X"53",X"95",X"B5",X"91",
		X"4E",X"3F",X"76",X"AD",X"A8",X"6A",X"3B",X"57",X"99",X"B3",X"8A",X"4A",X"41",X"7B",X"AF",X"A4",
		X"65",X"3A",X"5A",X"9B",X"B1",X"85",X"46",X"42",X"7E",X"AF",X"A1",X"61",X"3A",X"5E",X"9F",X"B1",
		X"82",X"44",X"45",X"82",X"B1",X"9F",X"5E",X"3A",X"61",X"A1",X"B0",X"7E",X"42",X"46",X"85",X"B2",
		X"9D",X"5C",X"3A",X"63",X"A2",X"B0",X"7D",X"41",X"46",X"85",X"B1",X"9B",X"5A",X"39",X"63",X"A2",
		X"AF",X"7C",X"41",X"47",X"85",X"B1",X"9B",X"59",X"39",X"63",X"A1",X"AE",X"7B",X"40",X"46",X"85",
		X"B0",X"9B",X"59",X"39",X"63",X"A1",X"AE",X"7C",X"40",X"46",X"84",X"B0",X"9B",X"59",X"38",X"62",
		X"A1",X"AE",X"7C",X"41",X"45",X"84",X"B0",X"9C",X"5B",X"39",X"61",X"A0",X"AF",X"7D",X"41",X"44",
		X"82",X"B0",X"9D",X"5C",X"38",X"5F",X"9F",X"AF",X"7F",X"42",X"43",X"80",X"AF",X"9E",X"5E",X"38",
		X"5C",X"9C",X"AF",X"81",X"43",X"41",X"7C",X"AE",X"A0",X"60",X"38",X"59",X"9A",X"B0",X"85",X"45",
		X"3F",X"79",X"AC",X"A2",X"63",X"37",X"55",X"96",X"B0",X"88",X"48",X"3D",X"74",X"AB",X"A5",X"69",
		X"39",X"51",X"92",X"B0",X"8C",X"4B",X"3A",X"6F",X"A8",X"A7",X"6E",X"3A",X"4D",X"8D",X"B1",X"92",
		X"50",X"39",X"69",X"A5",X"AA",X"73",X"3B",X"47",X"87",X"AF",X"96",X"54",X"37",X"63",X"A1",X"AC",
		X"79",X"3E",X"44",X"82",X"AF",X"9B",X"59",X"36",X"5C",X"9C",X"AE",X"7F",X"41",X"3F",X"7A",X"AC",
		X"A0",X"62",X"37",X"55",X"96",X"B0",X"88",X"47",X"3B",X"71",X"A8",X"A5",X"6A",X"38",X"4D",X"8E",
		X"B0",X"91",X"4F",X"38",X"68",X"A4",X"AB",X"74",X"3C",X"45",X"84",X"AE",X"98",X"57",X"36",X"5D",
		X"9C",X"AE",X"7F",X"42",X"3F",X"7A",X"AC",X"A1",X"62",X"36",X"53",X"93",X"AF",X"8A",X"49",X"39",
		X"6E",X"A7",X"A7",X"6E",X"3A",X"4A",X"8A",X"B0",X"94",X"53",X"37",X"62",X"A0",X"AC",X"7A",X"3E",
		X"41",X"7D",X"AD",X"9E",X"5F",X"36",X"56",X"96",X"AF",X"88",X"48",X"3B",X"70",X"A7",X"A6",X"6C",
		X"38",X"4A",X"8A",X"AF",X"93",X"52",X"36",X"62",X"A0",X"AC",X"7A",X"3E",X"41",X"7D",X"AD",X"9D",
		X"5E",X"35",X"55",X"95",X"AE",X"87",X"47",X"39",X"6F",X"A7",X"A6",X"6D",X"39",X"49",X"89",X"AF",
		X"94",X"53",X"35",X"5F",X"9D",X"AC",X"7D",X"40",X"3E",X"78",X"AB",X"A1",X"64",X"36",X"50",X"90",
		X"AF",X"8D",X"4C",X"37",X"67",X"A2",X"AA",X"75",X"3C",X"42",X"80",X"AD",X"9C",X"5D",X"35",X"56",
		X"97",X"AF",X"87",X"47",X"3A",X"6F",X"A7",X"A8",X"70",X"3A",X"48",X"88",X"B1",X"9A",X"59",X"38",
		X"5F",X"9E",X"B1",X"86",X"47",X"3F",X"77",X"AD",X"A9",X"6E",X"3C",X"4F",X"90",X"B5",X"99",X"58",
		X"3C",X"66",X"A4",X"B4",X"85",X"48",X"45",X"7F",X"B2",X"AA",X"6E",X"3F",X"56",X"96",X"B8",X"9A",
		X"59",X"40",X"6C",X"AA",X"B6",X"86",X"4A",X"4A",X"85",X"B6",X"AC",X"6F",X"42",X"5A",X"9B",X"BB",
		X"9C",X"5B",X"43",X"70",X"AD",X"B9",X"88",X"4C",X"4D",X"88",X"B9",X"AE",X"71",X"44",X"5D",X"9D",
		X"BD",X"9E",X"5D",X"45",X"72",X"AF",X"BB",X"8B",X"4F",X"4E",X"89",X"BB",X"B2",X"75",X"47",X"5E",
		X"9E",X"C0",X"A2",X"61",X"47",X"72",X"B0",X"BE",X"8F",X"52",X"4F",X"89",X"BD",X"B5",X"7A",X"49",
		X"5E",X"9E",X"C2",X"A7",X"66",X"48",X"71",X"AF",X"C1",X"94",X"56",X"4E",X"86",X"BC",X"B9",X"80",
		X"4C",X"5B",X"9A",X"C3",X"AC",X"6C",X"49",X"6C",X"AC",X"C3",X"9B",X"5C",X"4D",X"80",X"B9",X"BD",
		X"88",X"50",X"58",X"95",X"C2",X"B2",X"74",X"4A",X"67",X"A7",X"C4",X"A3",X"62",X"4C",X"7A",X"B6",
		X"C1",X"91",X"56",X"54",X"8D",X"C0",X"B9",X"7E",X"4D",X"61",X"A0",X"C5",X"AC",X"6C",X"4B",X"71",
		X"B0",X"C5",X"9C",X"5D",X"50",X"84",X"BD",X"C0",X"89",X"52",X"5A",X"97",X"C4",X"B5",X"76",X"4C",
		X"68",X"A8",X"C7",X"A6",X"66",X"4D",X"7A",X"B7",X"C4",X"95",X"58",X"54",X"8D",X"C1",X"BC",X"82",
		X"4F",X"5F",X"9E",X"C6",X"B0",X"71",X"4C",X"6E",X"AD",X"C7",X"A2",X"62",X"4F",X"7F",X"BA",X"C3",
		X"91",X"56",X"56",X"91",X"C3",X"BB",X"80",X"4F",X"62",X"A1",X"C8",X"AF",X"70",X"4D",X"71",X"B0",
		X"C8",X"A1",X"61",X"50",X"81",X"BB",X"C3",X"90",X"56",X"57",X"92",X"C3",X"BB",X"80",X"50",X"62",
		X"A1",X"C8",X"B0",X"71",X"4D",X"6F",X"AE",X"C7",X"A2",X"63",X"4F",X"7E",X"BA",X"C4",X"93",X"58",
		X"55",X"8E",X"C2",X"BD",X"84",X"51",X"5F",X"9D",X"C7",X"B4",X"75",X"4D",X"6B",X"AA",X"C8",X"A8",
		X"67",X"4E",X"78",X"B6",X"C6",X"9A",X"5D",X"52",X"87",X"BF",X"C1",X"8B",X"54",X"59",X"95",X"C5",
		X"B9",X"7D",X"4E",X"64",X"A3",X"C8",X"AF",X"6F",X"4D",X"70",X"AF",X"C8",X"A3",X"63",X"4E",X"7D",
		X"B9",X"C5",X"95",X"59",X"53",X"8A",X"C0",X"BF",X"87",X"52",X"5B",X"98",X"C5",X"B7",X"7A",X"4D",
		X"65",X"A4",X"C7",X"AC",X"6D",X"4C",X"70",X"AE",X"C6",X"A1",X"62",X"4E",X"7C",X"B7",X"C4",X"96",
		X"59",X"52",X"88",X"BE",X"BF",X"89",X"52",X"58",X"94",X"C3",X"B8",X"7D",X"4E",X"61",X"A0",X"C6",
		X"B0",X"71",X"4C",X"6C",X"AB",X"C7",X"A5",X"66",X"4C",X"76",X"B3",X"C5",X"9B",X"5C",X"4F",X"81",
		X"BB",X"C2",X"8F",X"55",X"54",X"8D",X"C0",X"BC",X"83",X"4F",X"5A",X"97",X"C4",X"B5",X"77",X"4B",
		X"62",X"A2",X"C6",X"AC",X"6D",X"4A",X"6C",X"AB",X"C6",X"A3",X"63",X"4B",X"76",X"B3",X"C4",X"99",
		X"5B",X"4E",X"80",X"B9",X"C1",X"8F",X"54",X"52",X"8B",X"BF",X"BC",X"84",X"4F",X"58",X"95",X"C2",
		X"B6",X"7A",X"4C",X"5F",X"9E",X"C4",X"AE",X"70",X"49",X"67",X"A6",X"C5",X"A6",X"67",X"4A",X"70",
		X"AE",X"C4",X"9E",X"5F",X"4B",X"78",X"B4",X"C2",X"95",X"58",X"4D",X"80",X"B9",X"BF",X"8C",X"53",
		X"51",X"89",X"BD",X"BB",X"84",X"4E",X"56",X"91",X"C0",X"B6",X"7A",X"4A",X"5B",X"99",X"C2",X"B0",
		X"72",X"48",X"62",X"A1",X"C3",X"AA",X"6A",X"48",X"69",X"A8",X"C3",X"A2",X"63",X"48",X"70",X"AD",
		X"C2",X"9B",X"5C",X"49",X"77",X"B3",X"C1",X"94",X"57",X"4C",X"7F",X"B7",X"BE",X"8C",X"51",X"4F",
		X"86",X"BB",X"BA",X"84",X"4D",X"53",X"8D",X"BE",X"B6",X"7C",X"4A",X"58",X"94",X"C0",X"B1",X"75",
		X"48",X"5C",X"9A",X"C1",X"AC",X"6E",X"46",X"61",X"A0",X"C1",X"A7",X"68",X"46",X"67",X"A5",X"C1",
		X"A1",X"62",X"46",X"6D",X"AA",X"C1",X"9B",X"5C",X"47",X"73",X"AF",X"BF",X"95",X"57",X"48",X"78",
		X"B3",X"BE",X"8F",X"53",X"4A",X"7E",X"B6",X"BB",X"89",X"4F",X"4C",X"83",X"B8",X"B8",X"83",X"4B",
		X"4E",X"88",X"BA",X"B5",X"7E",X"49",X"52",X"8D",X"BC",X"B2",X"78",X"47",X"55",X"92",X"BD",X"AF",
		X"72",X"45",X"58",X"96",X"BE",X"AB",X"6E",X"44",X"5C",X"9A",X"BF",X"A8",X"6A",X"43",X"60",X"9E",
		X"BF",X"A4",X"65",X"42",X"63",X"A1",X"BF",X"A0",X"61",X"42",X"67",X"A5",X"BE",X"9C",X"5D",X"43",
		X"6A",X"A7",X"BE",X"99",X"5A",X"43",X"6E",X"AA",X"BD",X"95",X"57",X"44",X"71",X"AC",X"BC",X"91",
		X"54",X"45",X"74",X"AE",X"BB",X"8E",X"52",X"45",X"77",X"B0",X"B9",X"8B",X"4F",X"46",X"79",X"B1",
		X"B8",X"88",X"4D",X"47",X"7C",X"B3",X"B8",X"86",X"4C",X"48",X"7E",X"B4",X"B6",X"83",X"4A",X"49",
		X"80",X"B5",X"B5",X"81",X"48",X"4A",X"82",X"B5",X"B4",X"7E",X"47",X"4B",X"84",X"B6",X"B3",X"7C",
		X"46",X"4B",X"85",X"B6",X"B1",X"7A",X"45",X"4C",X"86",X"B7",X"B1",X"79",X"45",X"4C",X"87",X"B7",
		X"B0",X"78",X"44",X"4D",X"87",X"B7",X"AF",X"77",X"43",X"4D",X"87",X"B6",X"AE",X"76",X"43",X"4D",
		X"88",X"B6",X"AE",X"76",X"43",X"4D",X"88",X"B6",X"AE",X"75",X"42",X"4D",X"88",X"B6",X"AD",X"74",
		X"42",X"4D",X"88",X"B6",X"AE",X"75",X"42",X"4C",X"87",X"B6",X"AE",X"75",X"42",X"4B",X"86",X"B5",
		X"AE",X"76",X"42",X"4A",X"85",X"B4",X"AE",X"77",X"43",X"4A",X"84",X"B4",X"AF",X"78",X"43",X"49",
		X"83",X"B4",X"AF",X"78",X"43",X"49",X"82",X"B4",X"B0",X"79",X"43",X"48",X"81",X"B3",X"B0",X"7A",
		X"44",X"47",X"80",X"B2",X"B1",X"7B",X"44",X"46",X"7E",X"B2",X"B2",X"7D",X"45",X"45",X"7C",X"B1",
		X"B2",X"7F",X"46",X"44",X"7A",X"B0",X"B3",X"81",X"47",X"43",X"78",X"AE",X"B4",X"83",X"49",X"42",
		X"76",X"AD",X"B5",X"86",X"4B",X"41",X"73",X"AB",X"B6",X"89",X"4D",X"40",X"6F",X"A9",X"B7",X"8C",
		X"4F",X"3F",X"6C",X"A7",X"B8",X"90",X"52",X"3E",X"68",X"A4",X"B8",X"94",X"55",X"3D",X"64",X"A1",
		X"B8",X"97",X"59",X"3C",X"60",X"9E",X"B9",X"9A",X"5C",X"3C",X"5D",X"9A",X"B9",X"9E",X"60",X"3C",
		X"59",X"97",X"B9",X"A1",X"64",X"3C",X"56",X"93",X"B8",X"A4",X"68",X"3D",X"52",X"8F",X"B7",X"A7",
		X"6C",X"3E",X"4F",X"8B",X"B6",X"AA",X"70",X"3F",X"4B",X"87",X"B5",X"AD",X"75",X"41",X"48",X"82",
		X"B3",X"B0",X"7A",X"44",X"45",X"7D",X"B0",X"B2",X"80",X"47",X"42",X"76",X"AD",X"B4",X"86",X"4B",
		X"40",X"71",X"AA",X"B6",X"8C",X"4F",X"3F",X"6B",X"A6",X"B7",X"91",X"53",X"3D",X"65",X"A1",X"B8",
		X"97",X"59",X"3C",X"5F",X"9C",X"B9",X"9C",X"5F",X"3C",X"5A",X"96",X"B8",X"A1",X"65",X"3D",X"54",
		X"90",X"B7",X"A6",X"6B",X"3E",X"4E",X"8A",X"B6",X"AB",X"73",X"41",X"4A",X"83",X"B3",X"B0",X"7A",
		X"44",X"45",X"7C",X"B0",X"B4",X"82",X"49",X"41",X"74",X"AC",X"B7",X"8B",X"4E",X"3E",X"6C",X"A6",
		X"B8",X"92",X"54",X"3C",X"64",X"A1",X"B9",X"99",X"5B",X"3C",X"5D",X"9A",X"BA",X"A0",X"63",X"3D",
		X"55",X"93",X"B8",X"A7",X"6B",X"3F",X"4E",X"8A",X"B6",X"AD",X"75",X"42",X"48",X"81",X"B2",X"B2",
		X"7F",X"47",X"43",X"77",X"AE",X"B6",X"88",X"4D",X"3F",X"6E",X"A8",X"B8",X"92",X"54",X"3D",X"64",
		X"A1",X"B9",X"9B",X"5D",X"3D",X"5B",X"98",X"B9",X"A3",X"66",X"3E",X"53",X"90",X"B8",X"AA",X"70",
		X"41",X"4B",X"86",X"B4",X"B0",X"7A",X"46",X"45",X"7C",X"AF",X"B5",X"85",X"4B",X"40",X"71",X"A9",
		X"B8",X"8F",X"53",X"3E",X"66",X"A2",X"BA",X"9A",X"5C",X"3D",X"5C",X"9A",X"B9",X"A4",X"66",X"3E",
		X"51",X"90",X"B7",X"AC",X"71",X"42",X"49",X"84",X"B3",X"B3",X"7E",X"47",X"43",X"78",X"AE",X"B7",
		X"89",X"4E",X"3F",X"6C",X"A7",X"B9",X"95",X"57",X"3D",X"61",X"9F",X"BA",X"A0",X"61",X"3E",X"56",
		X"95",X"B8",X"A9",X"6C",X"41",X"4C",X"89",X"B4",X"B1",X"79",X"46",X"45",X"7C",X"AF",X"B7",X"87",
		X"4D",X"40",X"6E",X"A8",X"B9",X"94",X"56",X"3E",X"61",X"9F",X"B9",X"A1",X"61",X"3F",X"55",X"94",
		X"B7",X"AB",X"6E",X"43",X"4A",X"87",X"B3",X"B3",X"7C",X"48",X"43",X"79",X"AE",X"B8",X"8B",X"50",
		X"40",X"6A",X"A6",X"B9",X"9A",X"5A",X"3F",X"5C",X"9C",X"B8",X"A6",X"66",X"41",X"4F",X"90",X"B5",
		X"B0",X"75",X"46",X"46",X"81",X"B1",X"B7",X"85",X"4C",X"41",X"70",X"AA",X"B9",X"95",X"55",X"3F",
		X"60",X"A1",X"B9",X"A4",X"61",X"41",X"52",X"95",X"B6",X"AF",X"70",X"45",X"48",X"85",X"B2",X"B6",
		X"81",X"4B",X"42",X"74",X"AC",X"B9",X"92",X"53",X"40",X"63",X"A4",X"B9",X"A2",X"5F",X"42",X"53",
		X"97",X"B6",X"AF",X"6E",X"46",X"48",X"87",X"B2",X"B6",X"80",X"4C",X"43",X"75",X"AC",X"B8",X"93",
		X"53",X"41",X"62",X"A4",X"B7",X"A4",X"5F",X"43",X"51",X"97",X"B4",X"B1",X"70",X"47",X"46",X"84",
		X"B1",X"B7",X"84",X"4D",X"42",X"70",X"AB",X"B8",X"98",X"55",X"42",X"5C",X"A1",X"B6",X"AA",X"63",
		X"45",X"4C",X"92",X"B3",X"B5",X"76",X"49",X"43",X"7D",X"AF",X"B9",X"8D",X"50",X"42",X"67",X"A8",
		X"B8",X"A1",X"5A",X"43",X"54",X"9D",X"B5",X"B0",X"6A",X"47",X"47",X"8A",X"B2",X"B8",X"80",X"4C",
		X"42",X"72",X"AD",X"B8",X"99",X"53",X"43",X"5A",X"A3",X"B5",X"AC",X"62",X"46",X"4A",X"92",X"B2",
		X"B7",X"78",X"4B",X"43",X"7A",X"AF",X"B8",X"91",X"50",X"43",X"61",X"A7",X"B5",X"A8",X"5D",X"47",
		X"4D",X"98",X"B2",X"B6",X"72",X"4A",X"44",X"80",X"AF",X"B8",X"8C",X"4F",X"43",X"65",X"AA",X"B5",
		X"A6",X"5A",X"47",X"4F",X"9C",X"B2",X"B6",X"6F",X"4B",X"44",X"83",X"AF",X"B9",X"8B",X"4F",X"43",
		X"66",X"AB",X"B5",X"A6",X"59",X"48",X"4E",X"9C",X"B1",X"B7",X"6F",X"4B",X"43",X"83",X"AF",X"B9",
		X"8C",X"4E",X"43",X"64",X"AB",X"B5",X"A8",X"5A",X"48",X"4C",X"9B",X"B1",X"B8",X"71",X"4B",X"43",
		X"80",X"B0",X"B9",X"90",X"4F",X"44",X"61",X"AA",X"B4",X"AB",X"5C",X"49",X"4A",X"99",X"B1",X"B9",
		X"75",X"4C",X"42",X"7B",X"AF",X"B9",X"95",X"51",X"46",X"5B",X"A8",X"B3",X"AF",X"60",X"4B",X"48",
		X"94",X"B0",X"BA",X"7C",X"4D",X"43",X"74",X"AF",X"B7",X"9C",X"53",X"48",X"55",X"A5",X"B1",X"B4",
		X"66",X"4C",X"44",X"8C",X"B0",X"BA",X"86",X"4E",X"44",X"69",X"AD",X"B5",X"A6",X"58",X"4A",X"4D",
		X"9E",X"B0",X"B8",X"70",X"4D",X"43",X"80",X"AF",X"B9",X"92",X"50",X"46",X"5D",X"AA",X"B3",X"B0",
		X"5F",X"4B",X"46",X"94",X"B0",X"BB",X"7E",X"4D",X"43",X"70",X"AE",X"B6",X"A1",X"54",X"48",X"50",
		X"A2",X"B1",X"B8",X"6B",X"4C",X"42",X"84",X"B0",X"BA",X"8F",X"4F",X"45",X"5E",X"AB",X"B3",X"AF",
		X"5D",X"4B",X"46",X"94",X"B0",X"BB",X"7E",X"4D",X"43",X"6F",X"AE",X"B6",X"A3",X"55",X"49",X"4E",
		X"A0",X"B0",X"B9",X"6F",X"4D",X"42",X"7F",X"AF",X"B9",X"95",X"50",X"47",X"59",X"A8",X"B1",X"B3",
		X"62",X"4C",X"44",X"8E",X"AF",X"BB",X"86",X"4E",X"44",X"66",X"AD",X"B4",X"AB",X"5A",X"4B",X"49",
		X"99",X"AF",X"BB",X"79",X"4E",X"43",X"73",X"AF",X"B7",X"A1",X"54",X"49",X"50",X"A2",X"B0",X"B9",
		X"6E",X"4E",X"42",X"80",X"AF",X"B9",X"96",X"51",X"47",X"58",X"A8",X"B1",X"B5",X"65",X"4D",X"43",
		X"8B",X"B0",X"BB",X"8B",X"4F",X"45",X"61",X"AC",X"B3",X"B0",X"5D",X"4C",X"45",X"93",X"B0",X"BC",
		X"82",X"4E",X"44",X"69",X"AE",X"B5",X"AA",X"59",X"4B",X"48",X"9A",X"B0",X"BC",X"7B",X"4D",X"43",
		X"70",X"AF",X"B6",X"A5",X"56",X"4A",X"4C",X"9F",X"B0",X"BB",X"75",X"4D",X"42",X"76",X"B0",X"B7",
		X"A0",X"54",X"49",X"4F",X"A1",X"B0",X"BA",X"71",X"4D",X"42",X"7B",X"B0",X"B8",X"9C",X"53",X"49",
		X"52",X"A4",X"B0",X"B9",X"6D",X"4D",X"42",X"7E",X"B0",X"B9",X"9A",X"52",X"49",X"54",X"A5",X"B0",
		X"B8",X"6B",X"4D",X"42",X"7F",X"B0",X"B9",X"99",X"52",X"48",X"54",X"A5",X"B0",X"B8",X"6C",X"4E",
		X"42",X"80",X"B0",X"B9",X"99",X"52",X"48",X"53",X"A5",X"B1",X"B9",X"6D",X"4E",X"42",X"7E",X"B0",
		X"B9",X"9B",X"52",X"48",X"52",X"A4",X"B1",X"B9",X"6D",X"4D",X"42",X"7D",X"B0",X"B9",X"9C",X"52",
		X"49",X"51",X"A3",X"B0",X"BA",X"70",X"4D",X"42",X"7A",X"B0",X"B8",X"9F",X"53",X"49",X"4E",X"A1",
		X"B0",X"BB",X"74",X"4D",X"42",X"75",X"B0",X"B7",X"A4",X"55",X"4A",X"4C",X"9E",X"B0",X"BB",X"79",
		X"4D",X"43",X"6F",X"AF",X"B6",X"A9",X"58",X"4B",X"48",X"99",X"B0",X"BC",X"80",X"4E",X"44",X"68",
		X"AE",X"B4",X"AE",X"5D",X"4C",X"45",X"91",X"B0",X"BC",X"89",X"4F",X"46",X"5F",X"AB",X"B2",X"B4",
		X"63",X"4D",X"43",X"88",X"B0",X"BB",X"93",X"50",X"47",X"56",X"A7",X"B1",X"B8",X"6B",X"4E",X"42",
		X"7E",X"B0",X"B8",X"9E",X"53",X"49",X"4F",X"A1",X"B0",X"BB",X"76",X"4D",X"42",X"71",X"AF",X"B6",
		X"A9",X"58",X"4B",X"48",X"97",X"B0",X"BC",X"83",X"4E",X"44",X"64",X"AD",X"B3",X"B2",X"60",X"4C",
		X"43",X"8B",X"B1",X"BB",X"92",X"50",X"47",X"57",X"A8",X"B1",X"B9",X"6C",X"4D",X"42",X"7B",X"B0",
		X"B8",X"A1",X"54",X"4A",X"4C",X"9E",X"B0",X"BC",X"7A",X"4D",X"43",X"6B",X"AF",X"B5",X"AD",X"5B",
		X"4C",X"45",X"91",X"B0",X"BC",X"8B",X"4F",X"46",X"5C",X"AA",X"B1",X"B7",X"68",X"4E",X"42",X"80",
		X"B0",X"B8",X"9E",X"53",X"4A",X"4D",X"9F",X"B0",X"BC",X"7B",X"4E",X"44",X"6A",X"AE",X"B4",X"AF",
		X"5D",X"4D",X"45",X"8E",X"B0",X"BB",X"90",X"50",X"47",X"57",X"A8",X"B1",X"B9",X"6D",X"4D",X"42",
		X"78",X"B0",X"B7",X"A5",X"56",X"4B",X"49",X"99",X"B0",X"BC",X"83",X"4E",X"45",X"61",X"AC",X"B3",
		X"B4",X"64",X"4D",X"42",X"84",X"B1",X"BA",X"9B",X"52",X"49",X"4E",X"A0",X"B1",X"BC",X"7A",X"4D",
		X"43",X"6A",X"AF",X"B5",X"B0",X"5E",X"4C",X"44",X"8B",X"B1",X"BB",X"94",X"50",X"48",X"53",X"A5",
		X"B1",X"BB",X"74",X"4D",X"43",X"70",X"B0",X"B5",X"AC",X"5B",X"4C",X"45",X"90",X"B0",X"BB",X"90",
		X"50",X"48",X"56",X"A7",X"B1",X"BA",X"71",X"4D",X"43",X"73",X"B0",X"B6",X"AA",X"5A",X"4C",X"46",
		X"91",X"B0",X"BB",X"8F",X"50",X"48",X"56",X"A7",X"B1",X"BA",X"71",X"4D",X"43",X"71",X"B0",X"B5",
		X"AC",X"5B",X"4C",X"45",X"8E",X"B0",X"BB",X"93",X"50",X"48",X"53",X"A4",X"B0",X"BB",X"76",X"4D",
		X"43",X"6D",X"AF",X"B4",X"AF",X"5E",X"4D",X"43",X"8A",X"B1",X"BB",X"98",X"51",X"49",X"4F",X"A1",
		X"B0",X"BC",X"7A",X"4D",X"43",X"68",X"AE",X"B4",X"B2",X"61",X"4D",X"42",X"85",X"B1",X"BA",X"9D",
		X"53",X"4A",X"4B",X"9D",X"B1",X"BD",X"82",X"4E",X"45",X"5F",X"AB",X"B2",X"B7",X"6A",X"4D",X"42",
		X"78",X"B1",X"B7",X"A8",X"58",X"4C",X"46",X"92",X"B1",X"BB",X"91",X"4F",X"48",X"53",X"A4",X"B1",
		X"BB",X"78",X"4D",X"44",X"69",X"AE",X"B3",X"B3",X"62",X"4D",X"43",X"82",X"B1",X"B9",X"A0",X"54",
		X"4B",X"4A",X"9A",X"B0",X"BC",X"88",X"4F",X"46",X"5A",X"A9",X"B1",X"B9",X"70",X"4E",X"43",X"71",
		X"B0",X"B5",X"AE",X"5D",X"4D",X"44",X"8A",X"B1",X"BA",X"9A",X"53",X"4A",X"4C",X"9D",X"B0",X"BD",
		X"84",X"4E",X"46",X"5D",X"AA",X"B2",X"B9",X"6E",X"4D",X"42",X"73",X"B0",X"B6",X"AE",X"5D",X"4D",
		X"43",X"89",X"B1",X"BA",X"9B",X"52",X"4A",X"4C",X"9D",X"B1",X"BD",X"84",X"4E",X"45",X"5D",X"AA",
		X"B2",X"B9",X"6E",X"4D",X"42",X"72",X"B0",X"B6",X"AE",X"5D",X"4C",X"43",X"88",X"B2",X"BA",X"9D",
		X"53",X"4A",X"4A",X"9A",X"B1",X"BD",X"89",X"4E",X"46",X"57",X"A7",X"B1",X"BB",X"75",X"4D",X"43",
		X"69",X"AF",X"B4",X"B4",X"64",X"4D",X"42",X"7C",X"B1",X"B7",X"A8",X"58",X"4C",X"45",X"8F",X"B1",
		X"BB",X"97",X"51",X"49",X"4D",X"9E",X"B0",X"BC",X"84",X"4E",X"46",X"5A",X"A9",X"B1",X"BA",X"72",
		X"4D",X"43",X"6C",X"AF",X"B3",X"B2",X"62",X"4D",X"42",X"7E",X"B1",X"B7",X"A6",X"57",X"4C",X"45",
		X"8F",X"B0",X"BB",X"97",X"51",X"49",X"4C",X"9D",X"B0",X"BC",X"86",X"4E",X"46",X"58",X"A8",X"B1",
		X"BB",X"75",X"4D",X"43",X"67",X"AE",X"B3",X"B6",X"67",X"4D",X"41",X"77",X"B1",X"B6",X"AD",X"5C",
		X"4C",X"42",X"86",X"B1",X"B9",X"A1",X"54",X"4B",X"46",X"94",X"B1",X"BC",X"93",X"4F",X"48",X"4E",
		X"A0",X"B1",X"BD",X"84",X"4D",X"46",X"58",X"A8",X"B1",X"BB",X"76",X"4D",X"43",X"65",X"AE",X"B3",
		X"B7",X"69",X"4D",X"42",X"73",X"B1",X"B5",X"AF",X"5F",X"4C",X"42",X"81",X"B1",X"B8",X"A6",X"57",
		X"4C",X"45",X"8E",X"B1",X"BA",X"9A",X"52",X"4A",X"4A",X"99",X"B1",X"BC",X"8E",X"4F",X"48",X"51",
		X"A2",X"B0",X"BC",X"82",X"4E",X"46",X"5A",X"A9",X"B1",X"BB",X"75",X"4D",X"43",X"65",X"AD",X"B2",
		X"B7",X"6A",X"4D",X"42",X"71",X"B0",X"B4",X"B2",X"61",X"4D",X"42",X"7D",X"B1",X"B7",X"AA",X"5A",
		X"4C",X"43",X"87",X"B1",X"B9",X"A2",X"55",X"4B",X"46",X"91",X"B1",X"BB",X"98",X"51",X"49",X"4A",
		X"9A",X"B1",X"BC",X"8E",X"4F",X"48",X"50",X"A1",X"B1",X"BD",X"84",X"4D",X"46",X"57",X"A7",X"B1",
		X"BC",X"7B",X"4C",X"44",X"5E",X"AB",X"B2",X"BA",X"72",X"4C",X"43",X"67",X"AE",X"B3",X"B7",X"6A",
		X"4C",X"42",X"6F",X"B0",X"B4",X"B3",X"63",X"4C",X"42",X"78",X"B1",X"B5",X"AE",X"5E",X"4C",X"42",
		X"80",X"B2",X"B7",X"A8",X"59",X"4C",X"43",X"88",X"B2",X"B9",X"A2",X"55",X"4B",X"45",X"8F",X"B1",
		X"BA",X"9B",X"52",X"4B",X"48",X"96",X"B1",X"BB",X"94",X"50",X"49",X"4C",X"9C",X"B1",X"BC",X"8C",
		X"4F",X"48",X"50",X"A1",X"B0",X"BD",X"86",X"4E",X"47",X"54",X"A4",X"B1",X"BD",X"81",X"4D",X"46",
		X"58",X"A7",X"B1",X"BC",X"7B",X"4D",X"45",X"5C",X"AA",X"B1",X"BB",X"77",X"4D",X"44",X"60",X"AC",
		X"B2",X"BA",X"73",X"4C",X"43",X"64",X"AD",X"B2",X"B9",X"6F",X"4C",X"43",X"67",X"AE",X"B3",X"B8",
		X"6C",X"4C",X"42",X"6B",X"AF",X"B3",X"B7",X"69",X"4C",X"42",X"6F",X"B0",X"B4",X"B5",X"66",X"4C",
		X"42",X"72",X"B1",X"B4",X"B3",X"64",X"4C",X"42",X"74",X"B1",X"B5",X"B2",X"62",X"4C",X"42",X"77",
		X"B1",X"B5",X"B1",X"61",X"4C",X"42",X"78",X"B1",X"B5",X"B0",X"60",X"4C",X"42",X"78",X"B1",X"B5",
		X"B0",X"60",X"4C",X"42",X"79",X"B1",X"B5",X"B0",X"60",X"4C",X"42",X"78",X"B1",X"B5",X"B0",X"60",
		X"4C",X"42",X"78",X"B1",X"B5",X"B1",X"61",X"4C",X"42",X"77",X"B1",X"B5",X"B1",X"61",X"4C",X"42",
		X"77",X"B1",X"B5",X"B1",X"61",X"4D",X"41",X"76",X"B1",X"B5",X"B2",X"62",X"4C",X"41",X"75",X"B1",
		X"B4",X"B3",X"63",X"4C",X"41",X"73",X"B1",X"B4",X"B4",X"65",X"4C",X"41",X"71",X"B0",X"B4",X"B5",
		X"66",X"4C",X"41",X"6F",X"B0",X"B4",X"B6",X"68",X"4C",X"42",X"6C",X"B0",X"B3",X"B7",X"6B",X"4C",
		X"42",X"69",X"AF",X"B3",X"B9",X"6E",X"4C",X"43",X"66",X"AE",X"B2",X"BA",X"71",X"4C",X"43",X"63",
		X"AD",X"B2",X"BB",X"74",X"4C",X"44",X"5F",X"AB",X"B2",X"BC",X"79",X"4C",X"45",X"5B",X"A9",X"B1",
		X"BC",X"7E",X"4C",X"46",X"56",X"A6",X"B1",X"BD",X"85",X"4D",X"47",X"52",X"A2",X"B1",X"BC",X"8A",
		X"4E",X"48",X"4E",X"9E",X"B1",X"BC",X"90",X"4F",X"49",X"4B",X"99",X"B1",X"BB",X"96",X"51",X"4A",
		X"48",X"94",X"B1",X"BA",X"9C",X"53",X"4B",X"45",X"8F",X"B2",X"B9",X"A2",X"55",X"4C",X"43",X"89",
		X"B2",X"B8",X"A7",X"59",X"4C",X"42",X"82",X"B2",X"B7",X"AD",X"5D",X"4C",X"41",X"7A",X"B1",X"B5",
		X"B2",X"63",X"4C",X"41",X"72",X"B0",X"B4",X"B6",X"69",X"4C",X"42",X"69",X"AF",X"B3",X"BA",X"71",
		X"4C",X"43",X"60",X"AC",X"B2",X"BC",X"7A",X"4C",X"45",X"57",X"A7",X"B1",X"BD",X"84",X"4D",X"47",
		X"50",X"A1",X"B1",X"BD",X"8F",X"4E",X"49",X"4A",X"99",X"B2",X"BB",X"99",X"51",X"4A",X"46",X"90",
		X"B2",X"B9",X"A3",X"56",X"4B",X"43",X"85",X"B2",X"B7",X"AB",X"5C",X"4C",X"42",X"79",X"B2",X"B4",
		X"B3",X"64",X"4C",X"42",X"6D",X"B0",X"B2",X"B8",X"6E",X"4C",X"43",X"62",X"AC",X"B1",X"BB",X"79",
		X"4C",X"45",X"58",X"A7",X"B1",X"BD",X"86",X"4E",X"48",X"4F",X"9E",X"B1",X"BC",X"93",X"50",X"4A",
		X"48",X"94",X"B2",X"BA",X"A0",X"55",X"4B",X"43",X"87",X"B2",X"B7",X"AB",X"5C",X"4C",X"41",X"79",
		X"B2",X"B5",X"B4",X"66",X"4C",X"42",X"6B",X"AF",X"B2",X"BA",X"72",X"4C",X"44",X"5D",X"AA",X"B1",
		X"BD",X"80",X"4C",X"46",X"51",X"A2",X"B1",X"BD",X"90",X"4F",X"49",X"48",X"96",X"B2",X"BB",X"9F",
		X"54",X"4B",X"43",X"88",X"B3",X"B8",X"AB",X"5C",X"4C",X"41",X"77",X"B2",X"B4",X"B5",X"68",X"4C",
		X"42",X"67",X"AE",X"B2",X"BB",X"76",X"4C",X"45",X"58",X"A7",X"B1",X"BD",X"88",X"4D",X"48",X"4C",
		X"9B",X"B2",X"BB",X"99",X"51",X"4B",X"45",X"8C",X"B3",X"B8",X"A9",X"5A",X"4C",X"42",X"7A",X"B2",
		X"B4",X"B4",X"66",X"4C",X"42",X"68",X"AE",X"B2",X"BB",X"76",X"4C",X"45",X"58",X"A6",X"B1",X"BD",
		X"88",X"4D",X"48",X"4B",X"9A",X"B1",X"BB",X"9B",X"53",X"4B",X"44",X"89",X"B2",X"B7",X"AB",X"5C",
		X"4C",X"41",X"76",X"B1",X"B4",X"B7",X"6B",X"4C",X"43",X"62",X"AC",X"B1",X"BC",X"7E",X"4C",X"46",
		X"51",X"A1",X"B1",X"BD",X"93",X"50",X"4A",X"46",X"90",X"B2",X"B9",X"A6",X"58",X"4C",X"41",X"7C",
		X"B2",X"B5",X"B4",X"66",X"4B",X"42",X"66",X"AE",X"B2",X"BC",X"7A",X"4C",X"46",X"54",X"A3",X"B2",
		X"BD",X"90",X"4E",X"49",X"47",X"92",X"B3",X"B9",X"A6",X"57",X"4B",X"41",X"7B",X"B2",X"B5",X"B5",
		X"68",X"4B",X"43",X"64",X"AD",X"B2",X"BC",X"7E",X"4C",X"47",X"51",X"A1",X"B2",X"BC",X"95",X"50",
		X"4A",X"45",X"8D",X"B3",X"B8",X"AA",X"5B",X"4C",X"42",X"75",X"B1",X"B3",X"B8",X"6E",X"4C",X"44",
		X"5D",X"AA",X"B1",X"BD",X"86",X"4D",X"49",X"4C",X"9A",X"B2",X"BB",X"9E",X"54",X"4C",X"43",X"83",
		X"B2",X"B6",X"B1",X"63",X"4C",X"42",X"69",X"AE",X"B2",X"BB",X"7A",X"4C",X"46",X"53",X"A2",X"B1",
		X"BD",X"94",X"50",X"4A",X"45",X"8C",X"B2",X"B8",X"AB",X"5C",X"4C",X"41",X"72",X"B1",X"B3",X"B9",
		X"71",X"4B",X"44",X"59",X"A7",X"B1",X"BD",X"8C",X"4E",X"49",X"47",X"93",X"B2",X"BA",X"A6",X"58",
		X"4B",X"41",X"79",X"B2",X"B4",X"B7",X"6B",X"4B",X"43",X"5D",X"AA",X"B2",X"BD",X"87",X"4D",X"48",
		X"4A",X"98",X"B2",X"BA",X"A2",X"55",X"4B",X"41",X"7D",X"B3",X"B5",X"B5",X"68",X"4B",X"43",X"60",
		X"AC",X"B1",X"BD",X"84",X"4C",X"48",X"4B",X"99",X"B2",X"BA",X"A0",X"55",X"4B",X"42",X"7E",X"B3",
		X"B4",X"B5",X"68",X"4C",X"43",X"60",X"AB",X"B1",X"BD",X"85",X"4D",X"49",X"4B",X"98",X"B2",X"BA",
		X"A2",X"56",X"4C",X"42",X"7A",X"B2",X"B4",X"B7",X"6C",X"4C",X"44",X"5C",X"A9",X"B1",X"BD",X"8A",
		X"4E",X"49",X"48",X"93",X"B3",X"B9",X"A7",X"5A",X"4C",X"41",X"74",X"B1",X"B3",X"B9",X"72",X"4C",
		X"45",X"57",X"A5",X"B1",X"BD",X"92",X"4F",X"4A",X"45",X"8B",X"B3",X"B7",X"AE",X"5F",X"4C",X"41",
		X"6B",X"AF",X"B2",X"BC",X"7B",X"4C",X"46",X"50",X"9F",X"B2",X"BC",X"9C",X"53",X"4B",X"42",X"81",
		X"B3",X"B5",X"B5",X"68",X"4B",X"42",X"5F",X"AB",X"B2",X"BD",X"88",X"4D",X"49",X"48",X"93",X"B3",
		X"B9",X"A8",X"5A",X"4B",X"41",X"71",X"B1",X"B3",X"BB",X"76",X"4B",X"46",X"52",X"A1",X"B2",X"BC",
		X"99",X"51",X"4B",X"42",X"82",X"B3",X"B5",X"B4",X"68",X"4B",X"43",X"5F",X"AA",X"B1",X"BD",X"8A",
		X"4D",X"49",X"47",X"91",X"B3",X"B8",X"AB",X"5D",X"4B",X"41",X"6B",X"AF",X"B2",X"BC",X"7D",X"4B",
		X"47",X"4D",X"9B",X"B2",X"BA",X"A2",X"56",X"4C",X"41",X"77",X"B2",X"B3",X"B9",X"72",X"4B",X"45",
		X"54",X"A3",X"B1",X"BC",X"98",X"51",X"4B",X"42",X"82",X"B3",X"B5",X"B5",X"69",X"4B",X"43",X"5C",
		X"A8",X"B1",X"BD",X"8F",X"4F",X"4A",X"44",X"8A",X"B3",X"B7",X"B1",X"63",X"4C",X"42",X"63",X"AC",
		X"B1",X"BD",X"88",X"4D",X"49",X"47",X"91",X"B3",X"B8",X"AC",X"5E",X"4C",X"41",X"69",X"AF",X"B2",
		X"BD",X"82",X"4C",X"48",X"49",X"96",X"B3",X"BA",X"A9",X"5B",X"4B",X"41",X"6C",X"B0",X"B2",X"BC",
		X"7F",X"4B",X"47",X"4B",X"98",X"B3",X"BA",X"A7",X"59",X"4B",X"41",X"6F",X"B1",X"B2",X"BC",X"7D",
		X"4B",X"47",X"4C",X"9A",X"B3",X"BA",X"A5",X"58",X"4B",X"41",X"71",X"B1",X"B2",X"BB",X"7B",X"4B",
		X"47",X"4D",X"9B",X"B2",X"BA",X"A4",X"58",X"4C",X"41",X"72",X"B1",X"B2",X"BB",X"7A",X"4B",X"47",
		X"4D",X"9B",X"B2",X"BA",X"A5",X"58",X"4C",X"41",X"71",X"B1",X"B2",X"BB",X"7B",X"4C",X"48",X"4C",
		X"99",X"B2",X"B9",X"A6",X"59",X"4C",X"41",X"6E",X"B0",X"B2",X"BC",X"7F",X"4C",X"48",X"4A",X"96",
		X"B3",X"B9",X"AA",X"5C",X"4B",X"41",X"69",X"AE",X"B2",X"BD",X"85",X"4C",X"48",X"47",X"91",X"B3",
		X"B8",X"AE",X"60",X"4B",X"42",X"63",X"AC",X"B1",X"BE",X"8A",X"4D",X"49",X"45",X"8C",X"B3",X"B7",
		X"B2",X"64",X"4B",X"42",X"5E",X"A9",X"B2",X"BD",X"91",X"4F",X"4A",X"43",X"85",X"B4",X"B5",X"B5",
		X"6A",X"4A",X"43",X"57",X"A6",X"B2",X"BD",X"99",X"51",X"4B",X"41",X"7D",X"B3",X"B4",X"B9",X"72",
		X"4A",X"45",X"51",X"A0",X"B3",X"BB",X"A1",X"56",X"4B",X"41",X"72",X"B1",X"B2",X"BC",X"7D",X"4B",
		X"48",X"4A",X"96",X"B3",X"B8",X"AB",X"5D",X"4B",X"42",X"66",X"AD",X"B2",X"BD",X"8A",X"4D",X"4A",
		X"45",X"8A",X"B3",X"B6",X"B3",X"67",X"4B",X"44",X"59",X"A7",X"B2",X"BC",X"99",X"52",X"4B",X"42",
		X"7A",X"B2",X"B3",X"BA",X"77",X"4B",X"47",X"4D",X"9A",X"B3",X"B9",X"A8",X"5A",X"4C",X"41",X"69",
		X"AE",X"B1",X"BD",X"88",X"4D",X"4A",X"45",X"8B",X"B3",X"B6",X"B3",X"67",X"4B",X"44",X"59",X"A6",
		X"B2",X"BD",X"9A",X"52",X"4B",X"41",X"78",X"B2",X"B3",X"BB",X"79",X"4B",X"47",X"4B",X"98",X"B3",
		X"B9",X"AB",X"5D",X"4B",X"41",X"64",X"AD",X"B2",X"BE",X"8E",X"4E",X"4A",X"43",X"84",X"B4",X"B5",
		X"B8",X"6E",X"4A",X"45",X"51",X"A0",X"B3",X"BB",X"A3",X"57",X"4B",X"41",X"6C",X"B0",X"B2",X"BD",
		X"86",X"4C",X"49",X"45",X"8B",X"B4",X"B6",X"B4",X"68",X"4A",X"44",X"57",X"A5",X"B2",X"BC",X"9D",
		X"53",X"4B",X"41",X"73",X"B1",X"B2",X"BC",X"80",X"4B",X"48",X"47",X"90",X"B4",X"B7",X"B1",X"64",
		X"4B",X"43",X"5A",X"A7",X"B2",X"BC",X"9A",X"52",X"4B",X"41",X"76",X"B2",X"B2",X"BC",X"7D",X"4B",
		X"48",X"48",X"92",X"B3",X"B7",X"B0",X"63",X"4B",X"43",X"5B",X"A7",X"B1",X"BC",X"9A",X"52",X"4C",
		X"41",X"75",X"B2",X"B2",X"BC",X"7F",X"4C",X"49",X"47",X"8F",X"B3",X"B6",X"B3",X"67",X"4B",X"44",
		X"56",X"A4",X"B2",X"BC",X"A0",X"55",X"4B",X"41",X"6D",X"B0",X"B2",X"BD",X"87",X"4D",X"4A",X"44",
		X"87",X"B4",X"B5",X"B7",X"6E",X"4A",X"45",X"50",X"9E",X"B3",X"BA",X"A7",X"5A",X"4B",X"41",X"66",
		X"AD",X"B2",X"BE",X"8F",X"4E",X"4A",X"42",X"7F",X"B4",X"B4",X"BA",X"76",X"4A",X"47",X"4B",X"97",
		X"B4",X"B9",X"AE",X"61",X"4B",X"43",X"5C",X"A8",X"B2",X"BD",X"9A",X"52",X"4B",X"41",X"73",X"B2",
		X"B2",X"BD",X"83",X"4C",X"49",X"45",X"8B",X"B4",X"B5",X"B6",X"6C",X"4A",X"45",X"51",X"9F",X"B3",
		X"BA",X"A7",X"5A",X"4B",X"41",X"64",X"AD",X"B2",X"BD",X"93",X"4F",X"4B",X"41",X"7A",X"B3",X"B2",
		X"BB",X"7D",X"4B",X"49",X"47",X"8F",X"B4",X"B6",X"B4",X"69",X"4A",X"45",X"52",X"A0",X"B2",X"BA",
		X"A7",X"5A",X"4B",X"42",X"63",X"AC",X"B1",X"BD",X"94",X"50",X"4B",X"41",X"77",X"B2",X"B2",X"BC",
		X"81",X"4C",X"49",X"45",X"8B",X"B4",X"B5",X"B6",X"6D",X"4A",X"46",X"4F",X"9C",X"B3",X"B9",X"AB",
		X"5E",X"4B",X"42",X"5D",X"A9",X"B2",X"BD",X"9B",X"53",X"4B",X"41",X"6F",X"B0",X"B2",X"BD",X"89",
		X"4D",X"4A",X"42",X"82",X"B4",X"B4",X"BB",X"77",X"4B",X"47",X"49",X"93",X"B4",X"B7",X"B3",X"67",
		X"4A",X"44",X"53",X"A1",X"B3",X"BB",X"A7",X"5A",X"4B",X"41",X"61",X"AB",X"B2",X"BD",X"98",X"51",
		X"4B",X"41",X"71",X"B2",X"B2",X"BD",X"88",X"4C",X"4A",X"43",X"82",X"B4",X"B4",X"BB",X"78",X"4A",
		X"48",X"48",X"91",X"B4",X"B6",X"B5",X"6A",X"4A",X"45",X"50",X"9D",X"B3",X"B9",X"AC",X"5F",X"4B",
		X"43",X"5B",X"A7",X"B2",X"BC",X"A0",X"56",X"4B",X"41",X"68",X"AE",X"B2",X"BD",X"93",X"50",X"4B",
		X"41",X"75",X"B2",X"B2",X"BD",X"86",X"4C",X"4A",X"43",X"83",X"B4",X"B3",X"BA",X"79",X"4B",X"48",
		X"47",X"8F",X"B4",X"B5",X"B6",X"6D",X"4A",X"46",X"4E",X"9A",X"B3",X"B8",X"AF",X"63",X"4B",X"44",
		X"56",X"A3",X"B2",X"BA",X"A6",X"5A",X"4B",X"42",X"5F",X"AA",X"B2",X"BD",X"9D",X"54",X"4B",X"40",
		X"69",X"AE",X"B1",X"BE",X"93",X"4F",X"4A",X"40",X"75",X"B2",X"B2",X"BD",X"87",X"4C",X"49",X"42",
		X"81",X"B4",X"B3",X"BB",X"7B",X"4B",X"48",X"46",X"8C",X"B4",X"B5",X"B8",X"70",X"4A",X"46",X"4A",
		X"95",X"B4",X"B7",X"B3",X"68",X"4A",X"45",X"50",X"9D",X"B4",X"B9",X"AD",X"60",X"4A",X"43",X"56",
		X"A4",X"B3",X"BB",X"A7",X"5B",X"4B",X"42",X"5E",X"A9",X"B2",X"BC",X"A0",X"55",X"4B",X"41",X"65",
		X"AD",X"B2",X"BD",X"99",X"52",X"4B",X"41",X"6C",X"B0",X"B2",X"BD",X"91",X"4F",X"4B",X"41",X"74",
		X"B2",X"B2",X"BD",X"89",X"4D",X"4A",X"42",X"7C",X"B3",X"B2",X"BC",X"83",X"4B",X"4A",X"43",X"82",
		X"B4",X"B3",X"BB",X"7C",X"4B",X"49",X"45",X"89",X"B4",X"B4",X"B9",X"76",X"4A",X"48",X"47",X"8E",
		X"B4",X"B5",X"B7",X"71",X"4A",X"47",X"49",X"93",X"B4",X"B6",X"B6",X"6D",X"4A",X"47",X"4C",X"96",
		X"B4",X"B7",X"B4",X"69",X"4A",X"46",X"4E",X"9A",X"B4",X"B8",X"B2",X"66",X"4A",X"45",X"50",X"9D",
		X"B3",X"B9",X"AF",X"62",X"4A",X"44",X"53",X"A0",X"B3",X"BA",X"AC",X"5F",X"4A",X"43",X"56",X"A3",
		X"B3",X"BA",X"AA",X"5D",X"4A",X"42",X"58",X"A5",X"B3",X"BB",X"A8",X"5B",X"4A",X"42",X"5A",X"A6",
		X"B3",X"BB",X"A6",X"5A",X"4A",X"41",X"5B",X"A7",X"B3",X"BB",X"A5",X"59",X"4A",X"42",X"5C",X"A8",
		X"B3",X"BB",X"A5",X"59",X"4A",X"42",X"5D",X"A8",X"B3",X"BB",X"A4",X"58",X"4A",X"42",X"5D",X"A8",
		X"B3",X"BB",X"A4",X"58",X"4A",X"42",X"5E",X"A8",X"B2",X"BB",X"A3",X"58",X"4B",X"42",X"5E",X"A9",
		X"B2",X"BB",X"A3",X"58",X"4B",X"42",X"5D",X"A8",X"B2",X"BB",X"A4",X"59",X"4B",X"42",X"5D",X"A8",
		X"B2",X"BB",X"A5",X"5A",X"4B",X"42",X"5B",X"A6",X"B2",X"BB",X"A7",X"5B",X"4B",X"43",X"59",X"A5",
		X"B2",X"BA",X"A9",X"5D",X"4B",X"43",X"57",X"A3",X"B3",X"BA",X"AB",X"5F",X"4A",X"44",X"54",X"A1",
		X"B3",X"B9",X"AE",X"62",X"4A",X"44",X"51",X"9E",X"B4",X"B8",X"B0",X"65",X"4A",X"45",X"4F",X"9B",
		X"B4",X"B8",X"B3",X"68",X"4A",X"45",X"4C",X"98",X"B4",X"B7",X"B5",X"6C",X"4A",X"46",X"4A",X"94",
		X"B5",X"B6",X"B7",X"6F",X"4A",X"47",X"48",X"91",X"B5",X"B6",X"B8",X"73",X"49",X"47",X"46",X"8C",
		X"B5",X"B5",X"BA",X"78",X"4A",X"48",X"44",X"87",X"B5",X"B4",X"BC",X"7D",X"4A",X"49",X"43",X"82",
		X"B5",X"B3",X"BD",X"83",X"4B",X"4A",X"42",X"7B",X"B4",X"B2",X"BD",X"8A",X"4C",X"4A",X"41",X"74",
		X"B2",X"B2",X"BE",X"91",X"4F",X"4B",X"41",X"6D",X"B0",X"B2",X"BD",X"98",X"51",X"4A",X"41",X"65",
		X"AD",X"B2",X"BC",X"A0",X"56",X"4B",X"42",X"5E",X"A8",X"B2",X"BA",X"A7",X"5B",X"4A",X"43",X"57",
		X"A3",X"B3",X"B9",X"AE",X"62",X"4A",X"45",X"4F",X"9B",X"B4",X"B7",X"B4",X"6A",X"4A",X"47",X"4A",
		X"93",X"B5",X"B5",X"B8",X"73",X"4A",X"48",X"46",X"8A",X"B4",X"B4",X"BB",X"7D",X"4B",X"49",X"43",
		X"80",X"B4",X"B2",X"BD",X"87",X"4C",X"4A",X"41",X"75",X"B2",X"B2",X"BE",X"93",X"50",X"4B",X"40",
		X"6A",X"AE",X"B2",X"BD",X"9D",X"54",X"4A",X"41",X"5F",X"A9",X"B3",X"BC",X"A7",X"5C",X"4A",X"43",
		X"55",X"A1",X"B4",X"B9",X"B0",X"64",X"49",X"45",X"4D",X"99",X"B5",X"B7",X"B6",X"6E",X"49",X"47",
		X"47",X"8D",X"B5",X"B4",X"BB",X"7B",X"4A",X"49",X"43",X"80",X"B4",X"B3",X"BD",X"89",X"4C",X"4A",
		X"41",X"72",X"B2",X"B2",X"BE",X"97",X"51",X"4B",X"41",X"64",X"AC",X"B2",X"BC",X"A3",X"58",X"4A",
		X"43",X"58",X"A4",X"B4",X"B9",X"AE",X"63",X"49",X"45",X"4D",X"98",X"B5",X"B6",X"B7",X"70",X"49",
		X"48",X"46",X"8A",X"B5",X"B3",X"BC",X"80",X"4B",X"4A",X"42",X"7A",X"B3",X"B2",X"BD",X"90",X"4F",
		X"4B",X"41",X"6A",X"AF",X"B2",X"BC",X"9F",X"56",X"4A",X"42",X"5B",X"A6",X"B3",X"BA",X"AC",X"61",
		X"4A",X"44",X"4E",X"99",X"B4",X"B6",X"B6",X"6F",X"49",X"48",X"46",X"89",X"B5",X"B3",X"BC",X"82",
		X"4B",X"4A",X"41",X"76",X"B2",X"B2",X"BE",X"94",X"50",X"4B",X"41",X"64",X"AC",X"B2",X"BC",X"A5",
		X"5A",X"4A",X"43",X"54",X"A0",X"B4",X"B8",X"B2",X"69",X"49",X"46",X"49",X"91",X"B5",X"B5",X"BB",
		X"7A",X"4A",X"49",X"42",X"7D",X"B4",X"B3",X"BE",X"8F",X"4E",X"4A",X"40",X"69",X"AE",X"B3",X"BD",
		X"A2",X"57",X"4A",X"42",X"57",X"A3",X"B4",X"B9",X"B1",X"66",X"49",X"46",X"4A",X"92",X"B5",X"B5",
		X"BA",X"79",X"49",X"49",X"42",X"7F",X"B5",X"B3",X"BE",X"8E",X"4D",X"4A",X"40",X"69",X"AE",X"B2",
		X"BC",X"A2",X"58",X"4A",X"43",X"56",X"A2",X"B4",X"B8",X"B2",X"69",X"49",X"47",X"48",X"8E",X"B6",
		X"B4",X"BC",X"7F",X"4A",X"4A",X"41",X"77",X"B3",X"B2",X"BD",X"96",X"51",X"4B",X"41",X"61",X"AA",
		X"B3",X"BA",X"AA",X"5F",X"4A",X"45",X"4F",X"99",X"B5",X"B6",X"B8",X"73",X"49",X"49",X"44",X"83",
		X"B5",X"B2",X"BD",X"8C",X"4D",X"4B",X"40",X"69",X"AE",X"B2",X"BC",X"A4",X"59",X"4A",X"43",X"54",
		X"9F",X"B4",X"B7",X"B4",X"6D",X"49",X"48",X"46",X"89",X"B5",X"B3",X"BD",X"86",X"4C",X"4B",X"40",
		X"6F",X"B0",X"B2",X"BD",X"9F",X"55",X"4A",X"42",X"57",X"A2",X"B4",X"B8",X"B2",X"69",X"49",X"47",
		X"47",X"8C",X"B5",X"B4",X"BD",X"83",X"4B",X"4A",X"40",X"71",X"B1",X"B3",X"BD",X"9E",X"55",X"4A",
		X"42",X"58",X"A3",X"B4",X"B9",X"B3",X"69",X"48",X"47",X"46",X"8C",X"B5",X"B4",X"BD",X"85",X"4B",
		X"4A",X"40",X"6F",X"B0",X"B3",X"BD",X"A0",X"56",X"4A",X"42",X"56",X"A1",X"B5",X"B8",X"B4",X"6C",
		X"48",X"48",X"45",X"89",X"B5",X"B3",X"BD",X"88",X"4C",X"4B",X"40",X"6B",X"AF",X"B3",X"BC",X"A4",
		X"5A",X"4A",X"44",X"51",X"9C",X"B5",X"B6",X"B7",X"73",X"49",X"49",X"42",X"7F",X"B4",X"B3",X"BD",
		X"93",X"50",X"4B",X"41",X"60",X"A9",X"B3",X"B9",X"AD",X"63",X"49",X"46",X"49",X"91",X"B5",X"B4",
		X"BB",X"81",X"4A",X"4B",X"40",X"71",X"B0",X"B2",X"BC",X"A0",X"57",X"4A",X"43",X"54",X"9F",X"B5",
		X"B7",X"B6",X"71",X"49",X"49",X"43",X"81",X"B4",X"B3",X"BD",X"92",X"4F",X"4B",X"41",X"60",X"A8",
		X"B3",X"BA",X"AE",X"64",X"49",X"46",X"48",X"8E",X"B5",X"B4",X"BC",X"85",X"4B",X"4B",X"40",X"6D",
		X"AE",X"B3",X"BC",X"A5",X"5B",X"4A",X"44",X"4F",X"9A",X"B5",X"B6",X"B9",X"79",X"49",X"4A",X"40",
		X"78",X"B2",X"B3",X"BD",X"9C",X"54",X"4A",X"41",X"57",X"A2",X"B5",X"B8",X"B5",X"6E",X"48",X"48",
		X"43",X"83",X"B4",X"B3",X"BD",X"92",X"4F",X"4B",X"40",X"5F",X"A8",X"B4",X"BA",X"B0",X"66",X"48",
		X"47",X"46",X"8B",X"B6",X"B4",X"BD",X"8C",X"4C",X"4B",X"40",X"65",X"AB",X"B4",X"BA",X"AD",X"62",
		X"48",X"46",X"48",X"8F",X"B6",X"B4",X"BC",X"87",X"4B",X"4B",X"40",X"69",X"AD",X"B3",X"BB",X"AA",
		X"5F",X"49",X"46",X"4A",X"93",X"B6",X"B4",X"BB",X"83",X"4A",X"4B",X"40",X"6C",X"AE",X"B3",X"BB",
		X"A8",X"5E",X"49",X"46",X"4B",X"94",X"B5",X"B4",X"BB",X"83",X"4A",X"4B",X"40",X"6D",X"AE",X"B3",
		X"BB",X"A8",X"5D",X"49",X"45",X"4C",X"94",X"B5",X"B4",X"BB",X"82",X"4A",X"4B",X"40",X"6D",X"AE",
		X"B3",X"BB",X"A8",X"5D",X"49",X"45",X"4B",X"93",X"B5",X"B4",X"BC",X"84",X"4A",X"4B",X"40",X"6B",
		X"AD",X"B3",X"BB",X"AA",X"5F",X"49",X"45",X"49",X"91",X"B5",X"B4",X"BC",X"87",X"4B",X"4B",X"3F",
		X"68",X"AC",X"B3",X"BB",X"AC",X"61",X"49",X"46",X"48",X"8E",X"B5",X"B4",X"BD",X"8A",X"4C",X"4B",
		X"3F",X"64",X"AA",X"B4",X"BA",X"AF",X"65",X"48",X"47",X"45",X"89",X"B5",X"B4",X"BD",X"90",X"4E",
		X"4B",X"40",X"5E",X"A7",X"B5",X"B9",X"B3",X"6C",X"47",X"48",X"42",X"81",X"B4",X"B4",X"BD",X"99",
		X"52",X"4A",X"41",X"55",X"A0",X"B5",X"B7",X"B8",X"76",X"47",X"4A",X"40",X"76",X"B2",X"B3",X"BC",
		X"A3",X"58",X"49",X"44",X"4E",X"97",X"B6",X"B5",X"BB",X"82",X"4A",X"4B",X"40",X"6B",X"AE",X"B4",
		X"BB",X"AB",X"61",X"48",X"47",X"47",X"8D",X"B5",X"B3",X"BC",X"8E",X"4D",X"4B",X"41",X"5F",X"A7",
		X"B4",X"B8",X"B3",X"6D",X"48",X"49",X"42",X"7F",X"B3",X"B3",X"BD",X"9C",X"54",X"4B",X"43",X"52",
		X"9C",X"B5",X"B5",X"BA",X"7D",X"49",X"4B",X"40",X"6E",X"AE",X"B3",X"BB",X"AA",X"60",X"49",X"47",
		X"47",X"8D",X"B5",X"B3",X"BD",X"8F",X"4E",X"4B",X"40",X"5C",X"A5",X"B4",X"B8",X"B5",X"71",X"48",
		X"4A",X"41",X"79",X"B2",X"B3",X"BD",X"A1",X"58",X"49",X"44",X"4D",X"96",X"B6",X"B5",X"BC",X"85",
		X"4B",X"4B",X"3F",X"64",X"AA",X"B4",X"BA",X"B1",X"69",X"48",X"48",X"42",X"81",X"B4",X"B3",X"BE",
		X"9B",X"54",X"4A",X"42",X"51",X"9B",X"B6",X"B6",X"BB",X"7F",X"49",X"4B",X"3F",X"6A",X"AD",X"B4",
		X"BB",X"AE",X"65",X"48",X"47",X"44",X"85",X"B5",X"B3",X"BD",X"98",X"52",X"4A",X"42",X"53",X"9D",
		X"B6",X"B6",X"BA",X"7E",X"49",X"4B",X"3F",X"6A",X"AD",X"B4",X"BA",X"AE",X"65",X"48",X"48",X"44",
		X"85",X"B5",X"B3",X"BD",X"99",X"52",X"4A",X"42",X"52",X"9C",X"B6",X"B5",X"BA",X"80",X"49",X"4B",
		X"3F",X"68",X"AC",X"B4",X"B9",X"B0",X"68",X"47",X"49",X"43",X"80",X"B4",X"B3",X"BD",X"9E",X"56",
		X"4A",X"44",X"4F",X"97",X"B6",X"B4",X"BC",X"86",X"4B",X"4B",X"40",X"62",X"A8",X"B4",X"B8",X"B4",
		X"6F",X"48",X"4A",X"41",X"78",X"B2",X"B3",X"BC",X"A5",X"5B",X"49",X"46",X"49",X"8F",X"B5",X"B3",
		X"BD",X"91",X"4F",X"4B",X"41",X"58",X"A1",X"B5",X"B6",X"B9",X"7B",X"49",X"4B",X"3F",X"6C",X"AD",
		X"B4",X"BA",X"AF",X"66",X"48",X"48",X"43",X"81",X"B4",X"B3",X"BD",X"9E",X"56",X"49",X"44",X"4D",
		X"96",X"B6",X"B5",X"BD",X"8A",X"4C",X"4B",X"40",X"5D",X"A5",X"B5",X"B8",X"B7",X"75",X"47",X"4A",
		X"3F",X"71",X"B0",X"B4",X"BB",X"AC",X"62",X"48",X"47",X"44",X"84",X"B5",X"B3",X"BD",X"9D",X"55",
		X"49",X"43",X"4D",X"96",X"B6",X"B5",X"BD",X"8B",X"4C",X"4B",X"40",X"5C",X"A4",X"B5",X"B7",X"B8",
		X"77",X"47",X"4A",X"3F",X"6D",X"AE",X"B4",X"BA",X"AF",X"67",X"47",X"48",X"42",X"7F",X"B4",X"B3",
		X"BD",X"A2",X"58",X"49",X"45",X"4A",X"90",X"B6",X"B4",X"BD",X"92",X"4F",X"4A",X"42",X"55",X"9E",
		X"B6",X"B5",X"BA",X"81",X"49",X"4B",X"40",X"63",X"A9",X"B5",X"B8",X"B5",X"71",X"47",X"4A",X"40",
		X"72",X"B0",X"B3",X"BB",X"AC",X"63",X"47",X"48",X"43",X"82",X"B4",X"B3",X"BC",X"A0",X"57",X"49",
		X"45",X"4A",X"90",X"B6",X"B3",X"BD",X"93",X"4F",X"4B",X"42",X"54",X"9D",X"B5",X"B5",X"BB",X"84",
		X"4A",X"4B",X"40",X"60",X"A7",X"B5",X"B8",X"B7",X"75",X"48",X"4B",X"3F",X"6E",X"AE",X"B3",X"BA",
		X"AF",X"68",X"48",X"49",X"41",X"7B",X"B3",X"B3",X"BC",X"A6",X"5D",X"48",X"46",X"46",X"88",X"B5",
		X"B3",X"BD",X"9C",X"55",X"4A",X"44",X"4C",X"93",X"B6",X"B4",X"BE",X"91",X"4E",X"4A",X"41",X"54",
		X"9D",X"B6",X"B5",X"BC",X"86",X"4A",X"4B",X"40",X"5D",X"A5",X"B6",X"B7",X"B9",X"7B",X"48",X"4A",
		X"3F",X"67",X"AB",X"B5",X"B9",X"B4",X"70",X"47",X"4A",X"3F",X"71",X"B0",X"B4",X"BB",X"AF",X"67",
		X"47",X"49",X"41",X"7B",X"B3",X"B4",X"BC",X"A8",X"5F",X"47",X"47",X"44",X"84",X"B5",X"B3",X"BD",
		X"A1",X"58",X"48",X"46",X"48",X"8C",X"B6",X"B3",X"BD",X"99",X"53",X"49",X"44",X"4D",X"94",X"B6",
		X"B4",X"BD",X"92",X"4F",X"4A",X"43",X"52",X"9A",X"B6",X"B4",X"BC",X"8B",X"4C",X"4B",X"41",X"57",
		X"A0",X"B6",X"B5",X"BB",X"84",X"4A",X"4B",X"40",X"5D",X"A5",X"B5",X"B6",X"B9",X"7C",X"49",X"4C",
		X"40",X"63",X"A9",X"B4",X"B7",X"B6",X"76",X"48",X"4B",X"3F",X"69",X"AC",X"B4",X"B8",X"B4",X"71",
		X"48",X"4B",X"3F",X"6D",X"AE",X"B4",X"B9",X"B2",X"6D",X"47",X"4A",X"40",X"72",X"B0",X"B3",X"BA",
		X"B0",X"69",X"47",X"49",X"40",X"76",X"B1",X"B3",X"BB",X"AD",X"65",X"47",X"49",X"41",X"7B",X"B3",
		X"B3",X"BC",X"AA",X"62",X"48",X"48",X"42",X"7E",X"B3",X"B3",X"BC",X"A7",X"5E",X"48",X"47",X"44",
		X"83",X"B4",X"B3",X"BD",X"A4",X"5B",X"48",X"46",X"45",X"86",X"B5",X"B4",X"BD",X"A1",X"59",X"48",
		X"45",X"46",X"89",X"B6",X"B3",X"BD",X"9F",X"57",X"48",X"45",X"47",X"8B",X"B6",X"B4",X"BE",X"9E",
		X"56",X"48",X"45",X"48",X"8C",X"B6",X"B4",X"BE",X"9D",X"55",X"48",X"45",X"49",X"8E",X"B6",X"B4",
		X"BD",X"9C",X"54",X"48",X"45",X"49",X"8E",X"B7",X"B4",X"BD",X"9B",X"54",X"49",X"45",X"49",X"8E",
		X"B6",X"B3",X"BD",X"9C",X"55",X"49",X"45",X"49",X"8D",X"B6",X"B3",X"BD",X"9C",X"55",X"49",X"45",
		X"49",X"8D",X"B6",X"B3",X"BD",X"9D",X"56",X"49",X"46",X"48",X"8C",X"B6",X"B3",X"BD",X"9E",X"57",
		X"49",X"46",X"47",X"8A",X"B6",X"B3",X"BD",X"A0",X"58",X"49",X"46",X"46",X"88",X"B5",X"B3",X"BD",
		X"A2",X"5A",X"48",X"47",X"45",X"85",X"B5",X"B3",X"BC",X"A5",X"5C",X"48",X"47",X"43",X"81",X"B4",
		X"B3",X"BC",X"A8",X"60",X"47",X"48",X"42",X"7D",X"B3",X"B3",X"BB",X"AB",X"64",X"47",X"49",X"41",
		X"78",X"B2",X"B4",X"BB",X"AF",X"68",X"47",X"4A",X"40",X"73",X"B0",X"B4",X"BA",X"B2",X"6D",X"47",
		X"4A",X"3F",X"6E",X"AE",X"B4",X"B9",X"B4",X"71",X"47",X"4A",X"3F",X"69",X"AC",X"B5",X"B8",X"B7",
		X"77",X"47",X"4B",X"3F",X"63",X"A9",X"B6",X"B7",X"B9",X"7D",X"48",X"4B",X"3F",X"5E",X"A5",X"B6",
		X"B7",X"BB",X"83",X"49",X"4A",X"40",X"58",X"A1",X"B7",X"B6",X"BC",X"8A",X"4B",X"4A",X"41",X"53",
		X"9B",X"B7",X"B5",X"BD",X"91",X"4F",X"49",X"43",X"4E",X"95",X"B7",X"B4",X"BE",X"98",X"53",X"49",
		X"44",X"49",X"8D",X"B7",X"B3",X"BD",X"A0",X"58",X"48",X"46",X"45",X"85",X"B5",X"B3",X"BC",X"A7",
		X"5F",X"47",X"48",X"42",X"7B",X"B3",X"B4",X"BB",X"AE",X"67",X"47",X"4A",X"40",X"71",X"B0",X"B4",
		X"B9",X"B3",X"70",X"47",X"4B",X"3F",X"67",X"AB",X"B5",X"B7",X"B8",X"7B",X"48",X"4B",X"40",X"5E",
		X"A4",X"B6",X"B5",X"BB",X"86",X"4B",X"4B",X"41",X"54",X"9C",X"B6",X"B4",X"BD",X"92",X"50",X"4A",
		X"44",X"4C",X"92",X"B6",X"B3",X"BD",X"9D",X"56",X"49",X"46",X"45",X"86",X"B5",X"B3",X"BC",X"A8",
		X"60",X"47",X"48",X"41",X"78",X"B1",X"B3",X"BA",X"B1",X"6C",X"47",X"4A",X"3F",X"6A",X"AC",X"B5",
		X"B8",X"B8",X"7A",X"48",X"4B",X"3F",X"5D",X"A4",X"B6",X"B6",X"BC",X"88",X"4B",X"4A",X"41",X"51",
		X"99",X"B7",X"B4",X"BE",X"96",X"52",X"49",X"44",X"48",X"8C",X"B6",X"B3",X"BD",X"A3",X"5B",X"47",
		X"47",X"42",X"7E",X"B4",X"B4",X"BC",X"AE",X"67",X"46",X"49",X"3F",X"6F",X"AF",X"B5",X"B9",X"B6",
		X"75",X"47",X"4A",X"3F",X"61",X"A7",X"B6",X"B6",X"BB",X"85",X"4A",X"4A",X"41",X"53",X"9B",X"B7",
		X"B4",X"BD",X"95",X"51",X"49",X"44",X"49",X"8C",X"B7",X"B4",X"BD",X"A4",X"5C",X"47",X"48",X"42",
		X"7B",X"B3",X"B4",X"BB",X"B1",X"6C",X"46",X"4A",X"3F",X"68",X"AB",X"B6",X"B7",X"B9",X"7E",X"48",
		X"4B",X"40",X"57",X"9F",X"B7",X"B4",X"BD",X"92",X"4F",X"49",X"44",X"4A",X"8E",X"B7",X"B3",X"BD",
		X"A3",X"5B",X"47",X"48",X"42",X"7B",X"B3",X"B4",X"BA",X"B1",X"6D",X"47",X"4B",X"3F",X"67",X"AA",
		X"B5",X"B6",X"BA",X"81",X"4A",X"4B",X"41",X"54",X"9C",X"B7",X"B4",X"BD",X"96",X"52",X"49",X"45",
		X"47",X"88",X"B5",X"B3",X"BC",X"A9",X"61",X"47",X"49",X"40",X"73",X"AF",X"B4",X"B9",X"B5",X"75",
		X"47",X"4B",X"3F",X"5D",X"A3",X"B6",X"B5",X"BC",X"8C",X"4D",X"4A",X"43",X"4C",X"91",X"B6",X"B3",
		X"BD",X"A2",X"5B",X"47",X"48",X"41",X"7A",X"B2",X"B4",X"BA",X"B3",X"6F",X"46",X"4A",X"3F",X"63",
		X"A8",X"B6",X"B6",X"BC",X"87",X"4B",X"4A",X"41",X"4F",X"96",X"B7",X"B4",X"BE",X"9E",X"57",X"48",
		X"46",X"43",X"7F",X"B4",X"B4",X"BB",X"B0",X"6B",X"46",X"4A",X"3F",X"66",X"AA",X"B6",X"B7",X"BB",
		X"83",X"4A",X"4A",X"41",X"51",X"98",X"B8",X"B4",X"BE",X"9C",X"56",X"47",X"46",X"43",X"80",X"B4",
		X"B4",X"BB",X"B0",X"6B",X"46",X"4A",X"3F",X"65",X"A9",X"B6",X"B6",X"BB",X"86",X"4A",X"4A",X"42",
		X"4F",X"95",X"B8",X"B4",X"BD",X"A0",X"59",X"47",X"48",X"42",X"7B",X"B3",X"B4",X"BA",X"B3",X"70",
		X"46",X"4B",X"3F",X"60",X"A6",X"B6",X"B5",X"BC",X"8C",X"4D",X"4A",X"43",X"4B",X"90",X"B7",X"B3",
		X"BD",X"A5",X"5E",X"47",X"49",X"41",X"74",X"B0",X"B4",X"B8",X"B6",X"78",X"48",X"4B",X"40",X"58",
		X"9F",X"B7",X"B4",X"BD",X"96",X"52",X"49",X"46",X"46",X"84",X"B5",X"B3",X"BB",X"AE",X"69",X"46",
		X"4B",X"3F",X"66",X"A9",X"B5",X"B6",X"BB",X"87",X"4C",X"4B",X"43",X"4D",X"92",X"B7",X"B3",X"BD",
		X"A4",X"5D",X"47",X"49",X"40",X"73",X"B0",X"B5",X"B9",X"B8",X"7A",X"48",X"4B",X"40",X"55",X"9C",
		X"B7",X"B4",X"BE",X"9B",X"55",X"48",X"47",X"43",X"7D",X"B3",X"B4",X"BA",X"B3",X"71",X"46",X"4B",
		X"3F",X"5D",X"A3",X"B7",X"B5",X"BE",X"92",X"50",X"49",X"44",X"46",X"87",X"B6",X"B4",X"BC",X"AD",
		X"67",X"46",X"4A",X"3F",X"67",X"AA",X"B6",X"B7",X"BC",X"87",X"4B",X"4A",X"42",X"4C",X"91",X"B7",
		X"B4",X"BD",X"A6",X"5E",X"46",X"49",X"3F",X"70",X"AF",X"B6",X"B8",X"B9",X"7E",X"48",X"4A",X"41",
		X"52",X"98",X"B8",X"B4",X"BE",X"A0",X"59",X"46",X"48",X"41",X"76",X"B1",X"B5",X"B9",X"B7",X"79",
		X"47",X"4B",X"40",X"55",X"9C",X"B8",X"B4",X"BE",X"9D",X"57",X"47",X"48",X"42",X"79",X"B2",X"B5",
		X"B9",X"B6",X"78",X"47",X"4B",X"40",X"56",X"9C",X"B7",X"B4",X"BD",X"9D",X"57",X"47",X"48",X"42",
		X"78",X"B2",X"B4",X"B8",X"B6",X"79",X"47",X"4B",X"41",X"55",X"9B",X"B7",X"B3",X"BD",X"9E",X"58",
		X"47",X"48",X"41",X"78",X"B1",X"B4",X"B8",X"B7",X"79",X"48",X"4B",X"41",X"54",X"9B",X"B7",X"B3",
		X"BD",X"9F",X"59",X"47",X"48",X"41",X"76",X"B1",X"B4",X"B8",X"B8",X"7C",X"48",X"4B",X"41",X"52",
		X"98",X"B7",X"B3",X"BD",X"A2",X"5C",X"47",X"49",X"40",X"71",X"AF",X"B5",X"B8",X"BA",X"81",X"49",
		X"4A",X"41",X"4E",X"93",X"B7",X"B3",X"BD",X"A7",X"60",X"46",X"49",X"3F",X"6B",X"AC",X"B6",X"B7",
		X"BC",X"88",X"4C",X"4A",X"43",X"49",X"8C",X"B6",X"B3",X"BC",X"AD",X"68",X"46",X"4A",X"3E",X"62",
		X"A7",X"B7",X"B5",X"BD",X"92",X"50",X"48",X"45",X"44",X"82",X"B5",X"B4",X"BB",X"B3",X"72",X"46",
		X"4A",X"3F",X"58",X"9F",X"B8",X"B4",X"BE",X"9C",X"57",X"47",X"48",X"41",X"76",X"B1",X"B5",X"B9",
		X"B9",X"7E",X"48",X"4A",X"41",X"4F",X"94",X"B8",X"B4",X"BD",X"A7",X"61",X"45",X"4A",X"3F",X"68",
		X"AB",X"B7",X"B6",X"BC",X"8D",X"4D",X"48",X"45",X"47",X"86",X"B6",X"B4",X"BB",X"B1",X"6F",X"46",
		X"4B",X"3F",X"5A",X"A0",X"B8",X"B4",X"BE",X"9C",X"56",X"47",X"48",X"41",X"75",X"B1",X"B5",X"B8",
		X"B9",X"80",X"49",X"4A",X"42",X"4D",X"91",X"B7",X"B3",X"BC",X"AA",X"65",X"46",X"4B",X"3F",X"64",
		X"A7",X"B7",X"B5",X"BD",X"92",X"51",X"48",X"46",X"44",X"7E",X"B4",X"B4",X"B9",X"B6",X"78",X"47",
		X"4B",X"41",X"52",X"98",X"B7",X"B3",X"BD",X"A6",X"60",X"46",X"4A",X"3F",X"68",X"AA",X"B6",X"B5",
		X"BC",X"8E",X"4F",X"49",X"45",X"45",X"82",X"B4",X"B4",X"BA",X"B4",X"75",X"47",X"4B",X"40",X"54",
		X"9A",X"B7",X"B3",X"BE",X"A4",X"5D",X"46",X"49",X"3F",X"6A",X"AB",X"B6",X"B6",X"BD",X"8D",X"4E",
		X"49",X"45",X"45",X"83",X"B5",X"B4",X"BA",X"B5",X"75",X"46",X"4B",X"40",X"53",X"98",X"B8",X"B4",
		X"BE",X"A6",X"60",X"46",X"4A",X"3E",X"66",X"A9",X"B7",X"B6",X"BE",X"92",X"50",X"48",X"46",X"43",
		X"7C",X"B3",X"B5",X"B9",X"B8",X"7C",X"48",X"4A",X"41",X"4E",X"92",X"B8",X"B4",X"BD",X"AC",X"67",
		X"45",X"4A",X"3E",X"5F",X"A4",X"B8",X"B5",X"BE",X"9A",X"55",X"46",X"48",X"41",X"74",X"B0",X"B6",
		X"B7",X"BA",X"85",X"4A",X"49",X"43",X"48",X"89",X"B7",X"B4",X"BB",X"B2",X"70",X"45",X"4B",X"40",
		X"55",X"9B",X"B8",X"B4",X"BD",X"A5",X"5F",X"45",X"4A",X"3F",X"66",X"A9",X"B7",X"B5",X"BD",X"94",
		X"51",X"47",X"47",X"42",X"79",X"B2",X"B5",X"B8",X"B9",X"81",X"49",X"4A",X"43",X"4A",X"8C",X"B7",
		X"B3",X"BB",X"B0",X"6E",X"45",X"4B",X"40",X"57",X"9D",X"B8",X"B3",X"BD",X"A3",X"5E",X"46",X"4A",
		X"3F",X"67",X"A9",X"B7",X"B5",X"BD",X"93",X"51",X"48",X"47",X"42",X"78",X"B1",X"B5",X"B7",X"BA",
		X"83",X"4A",X"4A",X"44",X"48",X"89",X"B6",X"B3",X"BA",X"B3",X"73",X"47",X"4B",X"41",X"52",X"97",
		X"B7",X"B3",X"BD",X"AA",X"65",X"46",X"4B",X"3F",X"5E",X"A3",X"B7",X"B4",X"BE",X"9E",X"59",X"46",
		X"49",X"3F",X"6B",X"AB",X"B6",X"B5",X"BD",X"92",X"51",X"48",X"47",X"42",X"79",X"B2",X"B5",X"B8",
		X"BB",X"84",X"4A",X"49",X"44",X"47",X"86",X"B6",X"B4",X"BA",X"B5",X"76",X"46",X"4A",X"41",X"4F",
		X"93",X"B8",X"B4",X"BD",X"AE",X"6A",X"45",X"4B",X"3F",X"58",X"9E",X"B8",X"B4",X"BE",X"A4",X"5F",
		X"45",X"49",X"3E",X"63",X"A7",X"B8",X"B5",X"BE",X"9A",X"56",X"46",X"48",X"40",X"70",X"AE",X"B7",
		X"B7",X"BD",X"8E",X"4E",X"47",X"46",X"42",X"7B",X"B3",X"B5",X"B8",X"BA",X"83",X"4A",X"49",X"44",
		X"47",X"86",X"B6",X"B5",X"BA",X"B6",X"78",X"47",X"4A",X"41",X"4D",X"91",X"B8",X"B4",X"BC",X"B0",
		X"6D",X"45",X"4B",X"40",X"54",X"9A",X"B9",X"B4",X"BD",X"AA",X"65",X"45",X"4B",X"3F",X"5B",X"A0",
		X"B8",X"B3",X"BD",X"A3",X"5E",X"45",X"4A",X"3F",X"63",X"A6",X"B8",X"B4",X"BD",X"9C",X"58",X"46",
		X"49",X"40",X"6B",X"AB",X"B7",X"B5",X"BD",X"95",X"53",X"47",X"48",X"40",X"72",X"AF",X"B6",X"B6",
		X"BC",X"8E",X"4F",X"48",X"47",X"43",X"79",X"B2",X"B5",X"B7",X"BA",X"87",X"4B",X"49",X"45",X"45",
		X"80",X"B4",X"B4",X"B8",X"B8",X"80",X"49",X"4A",X"44",X"48",X"87",X"B6",X"B4",X"BA",X"B6",X"7A",
		X"48",X"4A",X"42",X"4A",X"8B",X"B6",X"B3",X"BA",X"B4",X"75",X"46",X"4B",X"41",X"4E",X"91",X"B7",
		X"B3",X"BC",X"B2",X"71",X"46",X"4B",X"40",X"50",X"94",X"B8",X"B3",X"BC",X"AF",X"6C",X"45",X"4B",
		X"3F",X"53",X"98",X"B8",X"B3",X"BD",X"AD",X"6A",X"45",X"4B",X"3F",X"55",X"9A",X"B8",X"B4",X"BD",
		X"AB",X"67",X"45",X"4A",X"3F",X"57",X"9C",X"B8",X"B4",X"BE",X"AA",X"65",X"45",X"4A",X"3F",X"59",
		X"9E",X"B9",X"B4",X"BE",X"A8",X"63",X"44",X"4A",X"3E",X"5A",X"9F",X"B8",X"B4",X"BE",X"A7",X"62",
		X"45",X"4A",X"3F",X"5C",X"A0",X"B9",X"B4",X"BE",X"A6",X"61",X"44",X"4A",X"3E",X"5C",X"A1",X"B8",
		X"B4",X"BE",X"A6",X"61",X"44",X"4A",X"3F",X"5D",X"A2",X"B9",X"B4",X"BE",X"A6",X"61",X"44",X"4A",
		X"3F",X"5C",X"A1",X"B9",X"B4",X"BD",X"A6",X"61",X"44",X"4A",X"3F",X"5C",X"A0",X"B9",X"B4",X"BD",
		X"A7",X"63",X"45",X"4B",X"3F",X"5A",X"9E",X"B9",X"B3",X"BD",X"A8",X"64",X"44",X"4B",X"3F",X"58",
		X"9D",X"B8",X"B3",X"BD",X"AB",X"67",X"45",X"4B",X"40",X"56",X"9A",X"B8",X"B3",X"BC",X"AC",X"69",
		X"45",X"4B",X"40",X"54",X"98",X"B8",X"B3",X"BC",X"AE",X"6C",X"45",X"4B",X"41",X"52",X"96",X"B8",
		X"B3",X"BB",X"B0",X"6F",X"46",X"4B",X"41",X"4F",X"92",X"B7",X"B3",X"BB",X"B2",X"72",X"46",X"4B",
		X"42",X"4D",X"8F",X"B7",X"B3",X"BB",X"B4",X"76",X"47",X"4B",X"42",X"4A",X"8B",X"B6",X"B4",X"BA",
		X"B6",X"7B",X"48",X"4A",X"43",X"47",X"86",X"B5",X"B4",X"B9",X"B9",X"81",X"4A",X"49",X"44",X"44",
		X"80",X"B4",X"B5",X"B8",X"BB",X"87",X"4C",X"48",X"46",X"42",X"7A",X"B2",X"B6",X"B7",X"BD",X"8D",
		X"4F",X"47",X"47",X"40",X"73",X"AF",X"B6",X"B6",X"BE",X"94",X"53",X"46",X"48",X"3F",X"6C",X"AB",
		X"B8",X"B5",X"BE",X"9B",X"57",X"45",X"49",X"3E",X"64",X"A7",X"B8",X"B4",X"BE",X"A2",X"5D",X"44",
		X"4A",X"3E",X"5D",X"A1",X"B9",X"B4",X"BE",X"A8",X"64",X"44",X"4A",X"3F",X"56",X"9B",X"B9",X"B4",
		X"BD",X"AE",X"6C",X"44",X"4A",X"40",X"50",X"93",X"B8",X"B4",X"BB",X"B3",X"75",X"46",X"4A",X"42",
		X"4A",X"8A",X"B7",X"B5",X"B9",X"B8",X"7E",X"48",X"49",X"44",X"45",X"80",X"B4",X"B6",X"B8",X"BB",
		X"89",X"4D",X"47",X"47",X"42",X"75",X"B0",X"B7",X"B6",X"BD",X"94",X"52",X"46",X"49",X"3F",X"69",
		X"AA",X"B8",X"B4",X"BE",X"9F",X"5B",X"45",X"4A",X"3F",X"5F",X"A2",X"B9",X"B3",X"BD",X"A9",X"65",
		X"44",X"4B",X"40",X"54",X"98",X"B8",X"B3",X"BB",X"B1",X"71",X"46",X"4B",X"42",X"4C",X"8C",X"B7",
		X"B3",X"B9",X"B7",X"7D",X"48",X"4A",X"45",X"45",X"80",X"B4",X"B5",X"B7",X"BB",X"8A",X"4E",X"48",
		X"48",X"41",X"72",X"AE",X"B7",X"B5",X"BE",X"99",X"56",X"46",X"4A",X"3E",X"63",X"A5",X"B8",X"B3",
		X"BD",X"A6",X"62",X"45",X"4B",X"3F",X"56",X"9A",X"B8",X"B3",X"BC",X"B1",X"71",X"46",X"4A",X"42",
		X"4A",X"8A",X"B6",X"B4",X"B9",X"B9",X"81",X"4A",X"49",X"45",X"43",X"7A",X"B2",X"B6",X"B7",X"BD",
		X"92",X"51",X"46",X"48",X"3F",X"6A",X"AA",X"B8",X"B4",X"BE",X"A1",X"5D",X"45",X"4A",X"3E",X"5A",
		X"9E",X"B9",X"B4",X"BD",X"AE",X"6C",X"45",X"4A",X"41",X"4D",X"8F",X"B7",X"B4",X"BA",X"B7",X"7C",
		X"48",X"48",X"44",X"44",X"7E",X"B3",X"B6",X"B7",X"BD",X"90",X"50",X"46",X"48",X"3F",X"6B",X"AB",
		X"B8",X"B5",X"BE",X"A1",X"5C",X"44",X"4A",X"3E",X"5A",X"9E",X"B9",X"B4",X"BD",X"AF",X"6D",X"45",
		X"4A",X"41",X"4C",X"8E",X"B8",X"B5",X"B9",X"B8",X"7F",X"49",X"48",X"45",X"42",X"7A",X"B2",X"B7",
		X"B6",X"BD",X"94",X"53",X"45",X"49",X"3F",X"65",X"A7",X"B8",X"B4",X"BD",X"A7",X"63",X"44",X"4A",
		X"40",X"52",X"96",X"B8",X"B4",X"BA",X"B5",X"78",X"47",X"49",X"45",X"45",X"80",X"B4",X"B6",X"B7",
		X"BC",X"8F",X"50",X"46",X"48",X"3F",X"69",X"A9",X"B8",X"B4",X"BD",X"A4",X"5F",X"45",X"4A",X"40",
		X"54",X"99",X"B8",X"B4",X"BA",X"B4",X"75",X"47",X"49",X"44",X"46",X"82",X"B4",X"B5",X"B6",X"BC",
		X"8E",X"4F",X"47",X"49",X"40",X"6A",X"AA",X"B7",X"B4",X"BD",X"A4",X"5F",X"45",X"4A",X"40",X"53",
		X"98",X"B7",X"B4",X"BA",X"B5",X"76",X"48",X"49",X"45",X"45",X"81",X"B3",X"B6",X"B6",X"BD",X"90",
		X"51",X"47",X"49",X"3F",X"66",X"A8",X"B7",X"B4",X"BD",X"A8",X"63",X"46",X"4A",X"41",X"4F",X"94",
		X"B6",X"B5",X"B9",X"B8",X"7D",X"4A",X"48",X"46",X"42",X"78",X"B1",X"B6",X"B6",X"BD",X"99",X"56",
		X"46",X"49",X"3F",X"5C",X"A2",X"B7",X"B5",X"BB",X"B1",X"6C",X"47",X"49",X"43",X"47",X"89",X"B5",
		X"B6",X"B7",X"BC",X"89",X"4E",X"47",X"47",X"40",X"6B",X"AC",X"B7",X"B6",X"BD",X"A6",X"5F",X"46",
		X"48",X"41",X"50",X"97",X"B7",X"B6",X"B9",X"B8",X"7B",X"49",X"47",X"46",X"42",X"79",X"B1",X"B7",
		X"B7",X"BD",X"9B",X"56",X"46",X"48",X"40",X"59",X"A1",X"B7",X"B7",X"BA",X"B3",X"6F",X"47",X"47",
		X"44",X"45",X"85",X"B4",X"B7",X"B7",X"BD",X"90",X"50",X"47",X"47",X"40",X"63",X"A9",X"B7",X"B7",
		X"BA",X"AD",X"65",X"47",X"47",X"44",X"49",X"8E",X"B5",X"B7",X"B7",X"BB",X"88",X"4D",X"47",X"47",
		X"41",X"6A",X"AC",X"B6",X"B7",X"BB",X"A9",X"5F",X"47",X"47",X"43",X"4C",X"94",X"B5",X"B7",X"B7",
		X"BA",X"81",X"4B",X"47",X"47",X"41",X"70",X"AF",X"B6",X"B6",X"BB",X"A5",X"5B",X"47",X"47",X"44",
		X"4F",X"98",X"B5",X"B7",X"B7",X"BA",X"7D",X"4B",X"47",X"47",X"42",X"72",X"B0",X"B6",X"B7",X"BB",
		X"A4",X"5A",X"48",X"47",X"44",X"4F",X"9A",X"B4",X"B7",X"B7",X"BA",X"7C",X"4B",X"47",X"47",X"42",
		X"73",X"B0",X"B5",X"B7",X"BB",X"A3",X"5A",X"48",X"47",X"44",X"4F",X"9A",X"B4",X"B7",X"B6",X"BA",
		X"7C",X"4B",X"47",X"47",X"41",X"72",X"B0",X"B5",X"B7",X"BB",X"A5",X"5B",X"49",X"46",X"44",X"4D",
		X"99",X"B4",X"B8",X"B6",X"BB",X"7F",X"4C",X"47",X"47",X"41",X"6E",X"AE",X"B5",X"B8",X"BA",X"A9",
		X"5D",X"49",X"46",X"45",X"4A",X"94",X"B4",X"B8",X"B6",X"BC",X"86",X"4D",X"47",X"46",X"41",X"67",
		X"AD",X"B4",X"B9",X"B9",X"AF",X"62",X"49",X"45",X"46",X"46",X"8D",X"B4",X"B8",X"B7",X"BD",X"8E",
		X"4E",X"48",X"45",X"41",X"5E",X"A9",X"B4",X"B9",X"B8",X"B4",X"69",X"4A",X"45",X"46",X"43",X"83",
		X"B3",X"B7",X"B8",X"BC",X"9A",X"52",X"49",X"45",X"44",X"53",X"A2",X"B4",X"BA",X"B6",X"BA",X"76",
		X"4A",X"45",X"46",X"41",X"73",X"B1",X"B5",X"B9",X"BA",X"A8",X"5A",X"49",X"44",X"46",X"4A",X"96",
		X"B4",X"B9",X"B6",X"BC",X"86",X"4C",X"47",X"46",X"42",X"63",X"AC",X"B4",X"B9",X"B7",X"B2",X"65",
		X"4A",X"45",X"47",X"44",X"86",X"B4",X"B7",X"B7",X"BB",X"98",X"51",X"49",X"45",X"44",X"53",X"A2",
		X"B3",X"BA",X"B5",X"BA",X"77",X"4B",X"46",X"47",X"42",X"71",X"B1",X"B4",X"B9",X"B8",X"AA",X"5C",
		X"4A",X"45",X"47",X"47",X"92",X"B3",X"B8",X"B5",X"BC",X"8D",X"4E",X"48",X"46",X"43",X"5C",X"A9",
		X"B3",X"BA",X"B5",X"B7",X"6E",X"4B",X"46",X"48",X"42",X"7B",X"B2",X"B5",X"B7",X"BA",X"A3",X"57",
		X"4A",X"45",X"46",X"4B",X"99",X"B2",X"B8",X"B5",X"BC",X"85",X"4D",X"48",X"47",X"42",X"62",X"AC",
		X"B3",X"BA",X"B6",X"B5",X"68",X"4B",X"45",X"48",X"42",X"80",X"B2",X"B6",X"B7",X"BB",X"A1",X"55",
		X"4A",X"44",X"46",X"4B",X"9A",X"B2",X"B9",X"B5",X"BD",X"86",X"4D",X"48",X"46",X"42",X"60",X"AB",
		X"B3",X"BA",X"B6",X"B6",X"6A",X"4B",X"45",X"47",X"41",X"7C",X"B2",X"B5",X"B8",X"BA",X"A5",X"57",
		X"4A",X"44",X"46",X"49",X"97",X"B3",X"B9",X"B6",X"BD",X"8B",X"4E",X"48",X"45",X"42",X"5A",X"A8",
		X"B3",X"BB",X"B6",X"BA",X"72",X"4B",X"45",X"47",X"40",X"72",X"B1",X"B5",X"BA",X"B9",X"AD",X"5E",
		X"4B",X"43",X"47",X"44",X"8C",X"B3",X"B8",X"B7",X"BC",X"98",X"51",X"49",X"44",X"45",X"50",X"A0",
		X"B3",X"BB",X"B5",X"BC",X"80",X"4C",X"46",X"46",X"42",X"64",X"AD",X"B3",X"BB",X"B6",X"B6",X"6A",
		X"4A",X"44",X"47",X"41",X"79",X"B2",X"B5",X"B9",X"B9",X"A9",X"5A",X"4A",X"43",X"47",X"46",X"90",
		X"B3",X"B8",X"B6",X"BC",X"96",X"50",X"49",X"44",X"45",X"51",X"A1",X"B3",X"BA",X"B4",X"BC",X"81",
		X"4C",X"47",X"46",X"43",X"60",X"AC",X"B3",X"BB",X"B5",X"B8",X"6F",X"4B",X"45",X"48",X"42",X"73",
		X"B1",X"B4",X"B9",X"B7",X"AE",X"5F",X"4B",X"44",X"48",X"43",X"86",X"B3",X"B6",X"B7",X"BA",X"A0",
		X"55",X"4A",X"44",X"47",X"4A",X"97",X"B3",X"B9",X"B5",X"BD",X"90",X"4F",X"49",X"45",X"45",X"54",
		X"A3",X"B2",X"BA",X"B4",X"BC",X"7E",X"4C",X"47",X"47",X"42",X"61",X"AB",X"B2",X"BA",X"B5",X"B8",
		X"6F",X"4B",X"46",X"48",X"41",X"71",X"B0",X"B4",X"B9",X"B7",X"B1",X"63",X"4B",X"44",X"48",X"42",
		X"7F",X"B2",X"B5",X"B8",X"B9",X"A7",X"59",X"4B",X"44",X"47",X"45",X"8D",X"B3",X"B7",X"B7",X"BC",
		X"9D",X"53",X"4A",X"44",X"46",X"4A",X"98",X"B3",X"B9",X"B5",X"BD",X"90",X"4F",X"49",X"44",X"44",
		X"51",X"A1",X"B2",X"BA",X"B5",X"BD",X"84",X"4C",X"48",X"45",X"43",X"5B",X"A8",X"B3",X"BB",X"B5",
		X"BC",X"78",X"4C",X"46",X"46",X"41",X"65",X"AD",X"B3",X"BB",X"B6",X"B8",X"6D",X"4A",X"45",X"47",
		X"40",X"70",X"B0",X"B4",X"BA",X"B8",X"B3",X"64",X"4A",X"44",X"47",X"41",X"7B",X"B2",X"B5",X"B9",
		X"B9",X"AD",X"5E",X"4A",X"43",X"47",X"42",X"83",X"B3",X"B6",X"B8",X"BA",X"A6",X"58",X"4A",X"43",
		X"47",X"45",X"8C",X"B4",X"B8",X"B7",X"BB",X"A0",X"54",X"4A",X"43",X"47",X"48",X"93",X"B4",X"B9",
		X"B6",X"BC",X"98",X"50",X"49",X"44",X"46",X"4B",X"9A",X"B3",X"B9",X"B5",X"BD",X"90",X"4E",X"49",
		X"44",X"45",X"50",X"A0",X"B3",X"BA",X"B5",X"BD",X"89",X"4D",X"48",X"45",X"44",X"54",X"A4",X"B3",
		X"BA",X"B4",X"BC",X"83",X"4C",X"48",X"45",X"44",X"59",X"A7",X"B3",X"BB",X"B5",X"BC",X"7F",X"4C",
		X"47",X"46",X"43",X"5C",X"A9",X"B3",X"BA",X"B4",X"BB",X"7C",X"4B",X"47",X"46",X"43",X"5E",X"AA",
		X"B2",X"BA",X"B4",X"BB",X"79",X"4B",X"47",X"47",X"42",X"62",X"AC",X"B3",X"BA",X"B5",X"BA",X"75",
		X"4B",X"47",X"47",X"42",X"64",X"AD",X"B3",X"BA",X"B5",X"B9",X"73",X"4B",X"46",X"47",X"42",X"66",
		X"AD",X"B2",X"BA",X"B5",X"B9",X"72",X"4B",X"46",X"47",X"42",X"66",X"AD",X"B3",X"BA",X"B5",X"B9",
		X"72",X"4B",X"46",X"47",X"41",X"66",X"AD",X"B2",X"BA",X"B5",X"BA",X"73",X"4B",X"46",X"47",X"42",
		X"65",X"AD",X"B3",X"BB",X"B5",X"BA",X"74",X"4B",X"46",X"47",X"41",X"64",X"AC",X"B3",X"BB",X"B5",
		X"BA",X"75",X"4B",X"46",X"46",X"41",X"62",X"AC",X"B3",X"BB",X"B5",X"BB",X"78",X"4B",X"46",X"46",
		X"42",X"60",X"AB",X"B3",X"BB",X"B5",X"BC",X"7A",X"4B",X"47",X"46",X"42",X"5D",X"A9",X"B3",X"BB",
		X"B5",X"BC",X"7D",X"4B",X"47",X"45",X"43",X"5A",X"A8",X"B3",X"BB",X"B5",X"BD",X"82",X"4C",X"47",
		X"45",X"43",X"56",X"A5",X"B3",X"BB",X"B5",X"BD",X"87",X"4C",X"48",X"44",X"44",X"52",X"A1",X"B3",
		X"BA",X"B6",X"BD",X"8E",X"4E",X"48",X"44",X"45",X"4E",X"9C",X"B4",X"BA",X"B6",X"BD",X"94",X"4F",
		X"49",X"43",X"46",X"49",X"96",X"B4",X"B9",X"B6",X"BC",X"9B",X"52",X"49",X"43",X"47",X"46",X"90",
		X"B4",X"B8",X"B7",X"BB",X"A3",X"56",X"4A",X"43",X"48",X"44",X"87",X"B4",X"B6",X"B8",X"B9",X"AA",
		X"5C",X"4A",X"44",X"48",X"42",X"7D",X"B3",X"B5",X"B9",X"B7",X"B1",X"64",X"4A",X"45",X"48",X"41",
		X"72",X"B1",X"B4",X"BA",X"B6",X"B6",X"6D",X"4A",X"45",X"47",X"41",X"66",X"AD",X"B3",X"BA",X"B4",
		X"BA",X"78",X"4B",X"47",X"46",X"43",X"5C",X"A9",X"B3",X"BA",X"B4",X"BC",X"84",X"4C",X"48",X"45",
		X"45",X"52",X"A0",X"B3",X"B9",X"B4",X"BD",X"91",X"4F",X"49",X"44",X"47",X"4A",X"96",X"B3",X"B8",
		X"B6",X"BC",X"9F",X"55",X"4A",X"44",X"48",X"44",X"88",X"B3",X"B6",X"B8",X"B9",X"AB",X"5D",X"4B",
		X"44",X"48",X"41",X"78",X"B2",X"B4",X"BA",X"B6",X"B5",X"69",X"4B",X"46",X"47",X"41",X"69",X"AE",
		X"B3",X"BB",X"B5",X"BB",X"78",X"4B",X"47",X"46",X"42",X"5A",X"A7",X"B2",X"BA",X"B5",X"BD",X"88",
		X"4D",X"49",X"44",X"45",X"4E",X"9C",X"B3",X"B9",X"B6",X"BD",X"99",X"52",X"4A",X"43",X"47",X"45",
		X"8D",X"B3",X"B7",X"B8",X"BA",X"A8",X"5A",X"4A",X"43",X"47",X"41",X"7C",X"B2",X"B5",X"BA",X"B8",
		X"B4",X"67",X"4A",X"45",X"47",X"41",X"69",X"AF",X"B4",X"BB",X"B5",X"BB",X"79",X"4A",X"46",X"45",
		X"42",X"57",X"A6",X"B3",X"BB",X"B5",X"BE",X"8D",X"4E",X"49",X"43",X"46",X"4A",X"97",X"B4",X"B9",
		X"B7",X"BC",X"A1",X"55",X"49",X"43",X"47",X"42",X"83",X"B4",X"B6",X"B9",X"B8",X"B0",X"63",X"49",
		X"44",X"47",X"41",X"6D",X"B0",X"B4",X"BB",X"B5",X"BA",X"77",X"4A",X"46",X"46",X"43",X"58",X"A6",
		X"B3",X"BA",X"B5",X"BD",X"8D",X"4D",X"48",X"44",X"46",X"4A",X"96",X"B4",X"B8",X"B7",X"BB",X"A3",
		X"57",X"4A",X"43",X"48",X"43",X"7F",X"B4",X"B5",X"BA",X"B6",X"B3",X"68",X"4A",X"45",X"47",X"41",
		X"66",X"AD",X"B3",X"BB",X"B4",X"BC",X"80",X"4B",X"48",X"45",X"45",X"51",X"9F",X"B3",X"B9",X"B5",
		X"BC",X"99",X"52",X"4A",X"44",X"48",X"44",X"88",X"B4",X"B6",X"B8",X"B8",X"AE",X"61",X"4A",X"45",
		X"48",X"41",X"6D",X"B0",X"B3",X"BA",X"B4",X"BB",X"7A",X"4B",X"48",X"46",X"44",X"55",X"A2",X"B3",
		X"B9",X"B5",X"BC",X"95",X"50",X"4A",X"44",X"47",X"45",X"8B",X"B3",X"B6",X"B8",X"B9",X"AD",X"60",
		X"4A",X"45",X"48",X"41",X"6E",X"B0",X"B3",X"BA",X"B5",X"BB",X"79",X"4B",X"48",X"46",X"44",X"54",
		X"A2",X"B3",X"B9",X"B5",X"BD",X"96",X"51",X"4A",X"44",X"47",X"44",X"89",X"B3",X"B6",X"B9",X"B9",
		X"B0",X"62",X"4A",X"45",X"47",X"40",X"6A",X"AE",X"B3",X"BB",X"B5",X"BC",X"7F",X"4B",X"48",X"45",
		X"44",X"4F",X"9D",X"B3",X"B9",X"B6",X"BC",X"9E",X"54",X"4A",X"43",X"47",X"42",X"80",X"B3",X"B5",
		X"BA",X"B7",X"B5",X"6A",X"4A",X"45",X"46",X"41",X"60",X"AA",X"B3",X"BB",X"B5",X"BE",X"8B",X"4D",
		X"49",X"44",X"46",X"48",X"93",X"B4",X"B8",X"B8",X"BA",X"A9",X"5B",X"4A",X"43",X"47",X"40",X"72",
		X"B1",X"B4",X"BB",X"B6",X"BB",X"78",X"4A",X"47",X"45",X"44",X"53",X"A2",X"B4",X"BA",X"B6",X"BD",
		X"9B",X"52",X"49",X"43",X"47",X"42",X"82",X"B4",X"B5",X"BA",X"B7",X"B5",X"6A",X"49",X"45",X"46",
		X"42",X"5E",X"AA",X"B4",X"BB",X"B5",X"BD",X"8F",X"4E",X"49",X"43",X"47",X"46",X"8D",X"B5",X"B7",
		X"B9",X"B8",X"AF",X"62",X"49",X"44",X"47",X"41",X"67",X"AE",X"B3",X"BB",X"B5",X"BD",X"86",X"4C",
		X"48",X"44",X"46",X"4A",X"95",X"B5",X"B8",X"B7",X"B9",X"A9",X"5C",X"49",X"44",X"48",X"41",X"6E",
		X"B0",X"B3",X"BB",X"B4",X"BB",X"7E",X"4B",X"48",X"45",X"46",X"4D",X"9A",X"B4",X"B8",X"B6",X"BA",
		X"A5",X"59",X"4A",X"44",X"48",X"41",X"73",X"B2",X"B4",X"BA",X"B4",X"BA",X"7A",X"4A",X"48",X"45",
		X"45",X"4F",X"9D",X"B4",X"B8",X"B6",X"BB",X"A3",X"58",X"4A",X"44",X"48",X"41",X"75",X"B2",X"B3",
		X"BA",X"B5",X"BB",X"7A",X"4B",X"48",X"45",X"45",X"4F",X"9C",X"B3",X"B8",X"B6",X"BB",X"A4",X"59",
		X"4A",X"44",X"48",X"41",X"72",X"B1",X"B3",X"BA",X"B5",X"BC",X"7E",X"4C",X"48",X"45",X"45",X"4C",
		X"99",X"B3",X"B8",X"B7",X"BA",X"A8",X"5C",X"4A",X"44",X"48",X"40",X"6C",X"AF",X"B3",X"BB",X"B5",
		X"BD",X"84",X"4C",X"49",X"44",X"46",X"49",X"93",X"B4",X"B7",X"B8",X"B9",X"AE",X"61",X"4A",X"45",
		X"47",X"41",X"64",X"AC",X"B3",X"BB",X"B5",X"BE",X"8D",X"4E",X"49",X"43",X"47",X"45",X"8A",X"B4",
		X"B6",X"B9",X"B8",X"B4",X"69",X"4A",X"45",X"46",X"42",X"5B",X"A7",X"B3",X"BA",X"B5",X"BD",X"98",
		X"51",X"49",X"43",X"47",X"41",X"7E",X"B3",X"B5",X"BB",X"B6",X"BA",X"75",X"4A",X"47",X"45",X"44",
		X"51",X"9E",X"B4",X"B9",X"B7",X"BB",X"A5",X"58",X"49",X"43",X"47",X"40",X"6F",X"B0",X"B4",X"BC",
		X"B5",X"BD",X"83",X"4B",X"48",X"43",X"46",X"48",X"91",X"B5",X"B7",X"B9",X"B9",X"B0",X"64",X"49",
		X"44",X"46",X"42",X"5F",X"AA",X"B4",X"BB",X"B5",X"BD",X"95",X"50",X"49",X"43",X"48",X"42",X"7F",
		X"B4",X"B5",X"BB",X"B6",X"B9",X"74",X"49",X"47",X"45",X"45",X"50",X"9E",X"B5",X"B9",X"B7",X"BA",
		X"A7",X"5A",X"49",X"44",X"48",X"41",X"6A",X"AF",X"B3",X"BB",X"B4",X"BD",X"8A",X"4D",X"49",X"43",
		X"47",X"45",X"88",X"B5",X"B5",X"BA",X"B6",X"B6",X"6E",X"49",X"46",X"46",X"44",X"54",X"A1",X"B4",
		X"B9",X"B6",X"BB",X"A4",X"58",X"4A",X"44",X"48",X"41",X"6C",X"AF",X"B3",X"BB",X"B4",X"BD",X"8A",
		X"4D",X"49",X"43",X"48",X"45",X"87",X"B4",X"B5",X"B9",X"B6",X"B7",X"70",X"4A",X"47",X"46",X"45",
		X"52",X"9F",X"B4",X"B8",X"B6",X"BA",X"A7",X"5B",X"4A",X"45",X"48",X"41",X"67",X"AE",X"B3",X"BA",
		X"B4",X"BD",X"90",X"4F",X"4A",X"44",X"48",X"43",X"81",X"B4",X"B4",X"BA",X"B5",X"BA",X"76",X"4A",
		X"48",X"45",X"45",X"4D",X"98",X"B4",X"B7",X"B7",X"B9",X"AD",X"61",X"4A",X"45",X"47",X"42",X"5F",
		X"A9",X"B3",X"BA",X"B5",X"BD",X"99",X"53",X"4A",X"44",X"48",X"41",X"77",X"B2",X"B3",X"BB",X"B5",
		X"BC",X"81",X"4C",X"49",X"44",X"46",X"46",X"8D",X"B4",X"B6",X"B9",X"B7",X"B5",X"6C",X"4A",X"46",
		X"45",X"43",X"53",X"A0",X"B4",X"B9",X"B7",X"BB",X"A8",X"5B",X"4A",X"44",X"47",X"41",X"65",X"AD",
		X"B3",X"BB",X"B5",X"BE",X"95",X"50",X"49",X"43",X"47",X"41",X"79",X"B3",X"B4",X"BB",X"B5",X"BD",
		X"81",X"4B",X"48",X"43",X"46",X"46",X"8D",X"B5",X"B6",X"BA",X"B7",X"B7",X"6F",X"49",X"46",X"45",
		X"44",X"4F",X"9C",X"B5",X"B8",X"B8",X"BA",X"AC",X"60",X"49",X"44",X"46",X"41",X"5C",X"A8",X"B4",
		X"BB",X"B6",X"BC",X"9F",X"55",X"49",X"43",X"48",X"41",X"6D",X"B0",X"B4",X"BC",X"B5",X"BE",X"8F",
		X"4E",X"49",X"43",X"48",X"42",X"7D",X"B4",X"B5",X"BB",X"B5",X"BB",X"7F",X"4A",X"47",X"43",X"46",
		X"46",X"8C",X"B5",X"B6",X"BA",X"B6",X"B7",X"71",X"49",X"46",X"45",X"45",X"4E",X"9A",X"B5",X"B8",
		X"B8",X"B9",X"B0",X"64",X"49",X"45",X"46",X"43",X"57",X"A4",X"B4",X"B9",X"B6",X"BA",X"A6",X"5A",
		X"49",X"44",X"47",X"41",X"62",X"AB",X"B3",X"BA",X"B5",X"BC",X"9A",X"53",X"49",X"43",X"48",X"41",
		X"6F",X"B1",X"B4",X"BB",X"B4",X"BD",X"8F",X"4E",X"49",X"43",X"48",X"42",X"7B",X"B3",X"B4",X"BB",
		X"B4",X"BC",X"83",X"4B",X"49",X"44",X"48",X"44",X"86",X"B4",X"B4",X"BA",X"B5",X"BA",X"79",X"4A",
		X"48",X"45",X"47",X"48",X"90",X"B5",X"B6",X"B9",X"B6",X"B7",X"70",X"4A",X"47",X"46",X"45",X"4D",
		X"98",X"B5",X"B7",X"B8",X"B8",X"B2",X"68",X"49",X"46",X"46",X"43",X"52",X"9E",X"B4",X"B8",X"B7",
		X"B9",X"AD",X"62",X"4A",X"46",X"47",X"43",X"57",X"A3",X"B4",X"B9",X"B7",X"BB",X"A9",X"5E",X"4A",
		X"45",X"47",X"42",X"5C",X"A7",X"B3",X"B9",X"B6",X"BB",X"A5",X"5A",X"4A",X"44",X"47",X"41",X"60",
		X"A9",X"B3",X"BA",X"B5",X"BC",X"A1",X"57",X"4A",X"44",X"48",X"41",X"64",X"AC",X"B3",X"BA",X"B5",
		X"BD",X"9F",X"55",X"4A",X"44",X"48",X"41",X"67",X"AD",X"B3",X"BB",X"B5",X"BD",X"9B",X"53",X"49",
		X"43",X"47",X"40",X"69",X"AE",X"B3",X"BB",X"B5",X"BD",X"99",X"52",X"49",X"43",X"48",X"40",X"6C",
		X"AF",X"B4",X"BB",X"B5",X"BE",X"97",X"51",X"49",X"43",X"47",X"40",X"6E",X"B0",X"B4",X"BC",X"B5",
		X"BE",X"95",X"50",X"49",X"42",X"47",X"40",X"6F",X"B1",X"B4",X"BC",X"B5",X"BE",X"93",X"50",X"49",
		X"42",X"48",X"41",X"71",X"B1",X"B4",X"BC",X"B5",X"BE",X"93",X"4F",X"49",X"43",X"48",X"41",X"72",
		X"B2",X"B4",X"BC",X"B5",X"BD",X"92",X"4F",X"49",X"43",X"48",X"41",X"71",X"B2",X"B4",X"BB",X"B5",
		X"BD",X"92",X"4F",X"49",X"43",X"48",X"41",X"71",X"B2",X"B4",X"BB",X"B5",X"BD",X"94",X"50",X"49",
		X"43",X"48",X"41",X"70",X"B1",X"B4",X"BB",X"B4",X"BD",X"95",X"51",X"49",X"43",X"48",X"41",X"6D",
		X"B0",X"B4",X"BB",X"B4",X"BC",X"99",X"52",X"49",X"43",X"48",X"41",X"69",X"AE",X"B4",X"BB",X"B5",
		X"BC",X"9D",X"55",X"49",X"44",X"48",X"42",X"64",X"AC",X"B4",X"BA",X"B5",X"BB",X"A2",X"58",X"49",
		X"44",X"48",X"42",X"5E",X"A9",X"B4",X"B9",X"B5",X"BA",X"A7",X"5B",X"49",X"45",X"47",X"43",X"59",
		X"A5",X"B4",X"B9",X"B7",X"BA",X"AC",X"61",X"49",X"45",X"47",X"44",X"54",X"A0",X"B5",X"B8",X"B7",
		X"B8",X"B0",X"66",X"49",X"46",X"46",X"44",X"4F",X"9A",X"B5",X"B7",X"B8",X"B7",X"B5",X"6C",X"49",
		X"47",X"45",X"46",X"4A",X"93",X"B5",X"B6",X"B9",X"B6",X"B9",X"75",X"4A",X"48",X"44",X"47",X"46",
		X"8B",X"B5",X"B4",X"BA",X"B5",X"BB",X"7F",X"4B",X"49",X"43",X"47",X"43",X"80",X"B3",X"B3",X"BB",
		X"B4",X"BD",X"89",X"4D",X"49",X"43",X"48",X"41",X"75",X"B2",X"B3",X"BB",X"B5",X"BE",X"95",X"51",
		X"4A",X"43",X"48",X"41",X"69",X"AE",X"B3",X"BB",X"B5",X"BD",X"A0",X"56",X"49",X"44",X"47",X"41",
		X"5E",X"A8",X"B4",X"BA",X"B7",X"BB",X"A9",X"5E",X"49",X"45",X"46",X"42",X"54",X"A1",X"B5",X"B8",
		X"B8",X"B9",X"B2",X"68",X"49",X"46",X"45",X"44",X"4C",X"96",X"B5",X"B7",X"BA",X"B7",X"B8",X"74",
		X"49",X"47",X"43",X"46",X"45",X"89",X"B5",X"B5",X"BB",X"B5",X"BC",X"82",X"4B",X"48",X"43",X"47",
		X"42",X"7A",X"B4",X"B4",X"BC",X"B5",X"BE",X"93",X"50",X"49",X"43",X"47",X"40",X"69",X"AF",X"B4",
		X"BB",X"B6",X"BC",X"A1",X"57",X"48",X"43",X"46",X"41",X"5A",X"A5",X"B5",X"B9",X"B8",X"B9",X"AF",
		X"63",X"48",X"45",X"45",X"45",X"4E",X"99",X"B6",X"B7",X"BA",X"B7",X"B8",X"74",X"49",X"47",X"43",
		X"47",X"45",X"88",X"B6",X"B5",X"BB",X"B4",X"BC",X"85",X"4B",X"48",X"43",X"48",X"41",X"74",X"B2",
		X"B4",X"BB",X"B5",X"BD",X"99",X"52",X"49",X"43",X"48",X"41",X"62",X"AB",X"B5",X"BA",X"B6",X"BA",
		X"AA",X"5F",X"49",X"45",X"46",X"44",X"51",X"9D",X"B5",X"B7",X"B9",X"B6",X"B6",X"70",X"48",X"47",
		X"44",X"47",X"46",X"88",X"B5",X"B4",X"BB",X"B4",X"BC",X"87",X"4C",X"49",X"43",X"49",X"41",X"71",
		X"B1",X"B4",X"BB",X"B4",X"BC",X"9E",X"56",X"49",X"44",X"48",X"42",X"5B",X"A5",X"B4",X"B8",X"B7",
		X"B8",X"B0",X"67",X"48",X"47",X"46",X"46",X"4A",X"92",X"B5",X"B5",X"BA",X"B5",X"BB",X"7F",X"4B",
		X"49",X"44",X"48",X"42",X"79",X"B3",X"B3",X"BB",X"B4",X"BD",X"98",X"53",X"4A",X"44",X"48",X"41",
		X"5F",X"A8",X"B3",X"B8",X"B6",X"B9",X"AE",X"63",X"49",X"46",X"46",X"45",X"4C",X"95",X"B5",X"B5",
		X"BA",X"B6",X"BB",X"7C",X"4B",X"49",X"44",X"48",X"42",X"7B",X"B3",X"B3",X"BB",X"B4",X"BD",X"97",
		X"52",X"49",X"44",X"47",X"41",X"5F",X"A8",X"B4",X"B9",X"B7",X"BA",X"AE",X"63",X"49",X"46",X"45",
		X"44",X"4B",X"94",X"B5",X"B6",X"BA",X"B6",X"BB",X"7D",X"4A",X"49",X"43",X"47",X"41",X"79",X"B3",
		X"B4",X"BB",X"B5",X"BE",X"9A",X"53",X"49",X"43",X"47",X"41",X"5C",X"A7",X"B4",X"B9",X"B8",X"B9",
		X"B1",X"67",X"48",X"46",X"44",X"45",X"48",X"8E",X"B6",X"B6",X"BB",X"B5",X"BD",X"86",X"4C",X"49",
		X"42",X"47",X"40",X"6E",X"B0",X"B4",X"BB",X"B6",X"BC",X"A4",X"5A",X"48",X"44",X"46",X"43",X"52",
		X"9E",X"B5",X"B8",X"BA",X"B7",X"B8",X"75",X"49",X"48",X"43",X"47",X"43",X"80",X"B5",X"B5",X"BC",
		X"B5",X"BD",X"95",X"50",X"48",X"42",X"47",X"41",X"5F",X"A8",X"B5",X"BA",X"B8",X"B9",X"B1",X"67",
		X"48",X"46",X"44",X"46",X"48",X"8D",X"B6",X"B5",X"BB",X"B5",X"BD",X"8A",X"4C",X"49",X"43",X"48",
		X"41",X"69",X"AE",X"B5",X"BA",X"B6",X"BB",X"A9",X"5E",X"48",X"45",X"45",X"45",X"4D",X"97",X"B6",
		X"B6",X"BA",X"B5",X"BA",X"7D",X"49",X"48",X"43",X"49",X"42",X"76",X"B3",X"B4",X"BB",X"B5",X"BC",
		X"A0",X"57",X"48",X"44",X"47",X"43",X"54",X"9F",X"B6",X"B7",X"B9",X"B6",X"B7",X"75",X"49",X"48",
		X"43",X"48",X"43",X"7C",X"B4",X"B4",X"BB",X"B4",X"BC",X"9C",X"54",X"49",X"44",X"48",X"43",X"57",
		X"A2",X"B5",X"B7",X"B8",X"B6",X"B6",X"72",X"48",X"48",X"43",X"48",X"43",X"7E",X"B4",X"B4",X"BB",
		X"B4",X"BD",X"9A",X"53",X"49",X"44",X"48",X"43",X"58",X"A2",X"B5",X"B7",X"B8",X"B7",X"B7",X"73",
		X"49",X"49",X"44",X"48",X"42",X"7D",X"B3",X"B3",X"BA",X"B4",X"BC",X"9C",X"54",X"49",X"45",X"48",
		X"43",X"55",X"A0",X"B5",X"B7",X"B8",X"B7",X"B8",X"76",X"49",X"49",X"44",X"49",X"42",X"79",X"B2",
		X"B3",X"BA",X"B5",X"BC",X"A1",X"58",X"49",X"45",X"47",X"43",X"51",X"9B",X"B5",X"B6",X"B9",X"B6",
		X"BA",X"7E",X"4A",X"49",X"43",X"48",X"40",X"70",X"B0",X"B4",X"BA",X"B6",X"BC",X"A9",X"5E",X"49",
		X"46",X"46",X"45",X"4B",X"93",X"B5",X"B5",X"BA",X"B5",X"BD",X"88",X"4C",X"4A",X"42",X"48",X"40",
		X"65",X"AB",X"B4",X"B9",X"B7",X"BA",X"B0",X"66",X"48",X"47",X"44",X"46",X"45",X"88",X"B5",X"B5",
		X"BB",X"B5",X"BE",X"95",X"50",X"49",X"43",X"47",X"41",X"5A",X"A4",X"B5",X"B8",X"B9",X"B8",X"B7",
		X"73",X"48",X"48",X"42",X"47",X"41",X"7A",X"B3",X"B4",X"BB",X"B6",X"BD",X"A1",X"57",X"48",X"44",
		X"46",X"43",X"50",X"9B",X"B6",X"B7",X"BB",X"B6",X"BC",X"81",X"4A",X"49",X"42",X"48",X"40",X"6B",
		X"AE",X"B5",X"BA",X"B7",X"BA",X"AD",X"63",X"47",X"46",X"43",X"46",X"45",X"89",X"B5",X"B5",X"BB",
		X"B5",X"BD",X"95",X"50",X"48",X"42",X"47",X"42",X"58",X"A3",X"B6",X"B8",X"BA",X"B7",X"B9",X"78",
		X"48",X"48",X"42",X"49",X"40",X"73",X"B2",X"B5",X"BB",X"B6",X"BA",X"A9",X"5E",X"47",X"45",X"44",
		X"45",X"48",X"8E",X"B6",X"B6",X"BB",X"B5",X"BD",X"91",X"4E",X"49",X"43",X"48",X"42",X"5B",X"A5",
		X"B6",X"B8",X"B9",X"B7",X"B8",X"76",X"48",X"49",X"42",X"49",X"41",X"73",X"B1",X"B5",X"BA",X"B6",
		X"BA",X"A9",X"5F",X"48",X"46",X"45",X"46",X"47",X"8D",X"B6",X"B5",X"BB",X"B5",X"BC",X"94",X"4F",
		X"49",X"43",X"48",X"43",X"58",X"A2",X"B6",X"B7",X"B9",X"B6",X"B9",X"7B",X"49",X"49",X"42",X"49",
		X"41",X"6D",X"AF",X"B5",X"B9",X"B6",X"B9",X"AE",X"65",X"48",X"47",X"44",X"48",X"44",X"84",X"B4",
		X"B4",X"BA",X"B4",X"BC",X"9D",X"55",X"49",X"45",X"47",X"44",X"4F",X"99",X"B6",X"B6",X"BA",X"B5",
		X"BC",X"89",X"4C",X"4A",X"43",X"49",X"41",X"61",X"A8",X"B5",X"B8",X"B7",X"B7",X"B6",X"73",X"48",
		X"49",X"43",X"49",X"40",X"74",X"B0",X"B4",X"B9",X"B6",X"BA",X"AC",X"62",X"48",X"47",X"44",X"47",
		X"45",X"86",X"B4",X"B4",X"BA",X"B5",X"BD",X"9D",X"55",X"4A",X"44",X"46",X"44",X"4E",X"98",X"B5",
		X"B6",X"BA",X"B5",X"BC",X"8B",X"4D",X"4A",X"42",X"48",X"40",X"5B",X"A4",X"B5",X"B7",X"B9",X"B7",
		X"B9",X"7B",X"49",X"4A",X"42",X"49",X"40",X"6A",X"AD",X"B5",X"BA",X"B8",X"BA",X"B3",X"6B",X"48",
		X"47",X"42",X"47",X"41",X"7B",X"B3",X"B4",X"BA",X"B6",X"BC",X"A8",X"5E",X"49",X"46",X"44",X"45",
		X"46",X"8B",X"B5",X"B5",X"BB",X"B5",X"BD",X"9B",X"53",X"49",X"44",X"46",X"43",X"4E",X"98",X"B6",
		X"B6",X"BB",X"B6",X"BD",X"8E",X"4D",X"49",X"42",X"47",X"41",X"58",X"A2",X"B6",X"B8",X"BA",X"B7",
		X"BB",X"81",X"4A",X"49",X"41",X"48",X"40",X"63",X"A9",X"B5",X"B9",X"B9",X"B8",X"B7",X"75",X"47",
		X"48",X"41",X"48",X"3F",X"6D",X"AF",X"B5",X"BA",X"B8",X"BA",X"B2",X"6A",X"47",X"47",X"42",X"48",
		X"41",X"79",X"B3",X"B5",X"BB",X"B7",X"BC",X"AB",X"61",X"48",X"46",X"44",X"47",X"44",X"84",X"B5",
		X"B5",X"BB",X"B5",X"BC",X"A3",X"59",X"47",X"45",X"45",X"45",X"48",X"8E",X"B6",X"B6",X"BB",X"B5",
		X"BD",X"95",X"50",X"48",X"43",X"47",X"42",X"54",X"9E",X"B6",X"B7",X"BA",X"B6",X"BC",X"87",X"4B",
		X"49",X"42",X"49",X"41",X"5C",X"A5",X"B6",X"B8",X"B9",X"B6",X"B9",X"7F",X"49",X"49",X"42",X"49",
		X"40",X"62",X"A9",X"B6",X"B9",X"B8",X"B6",X"B7",X"78",X"47",X"49",X"42",X"49",X"40",X"68",X"AC",
		X"B5",X"B9",X"B8",X"B7",X"B5",X"72",X"47",X"49",X"42",X"4A",X"41",X"6F",X"AF",X"B5",X"B9",X"B7",
		X"B8",X"B3",X"6D",X"47",X"48",X"42",X"49",X"41",X"74",X"B1",X"B5",X"B9",X"B6",X"B8",X"B0",X"69",
		X"47",X"48",X"43",X"49",X"41",X"77",X"B2",X"B4",X"BA",X"B6",X"B9",X"AE",X"66",X"47",X"48",X"44",
		X"49",X"42",X"7A",X"B2",X"B4",X"B9",X"B6",X"BA",X"AD",X"64",X"47",X"48",X"44",X"49",X"42",X"7C",
		X"B3",X"B4",X"BA",X"B6",X"BA",X"AC",X"63",X"48",X"48",X"44",X"48",X"43",X"7E",X"B3",X"B4",X"BA",
		X"B5",X"BA",X"AB",X"61",X"48",X"48",X"44",X"48",X"42",X"7E",X"B3",X"B4",X"BA",X"B5",X"BB",X"AA",
		X"61",X"48",X"47",X"44",X"48",X"42",X"7E",X"B3",X"B4",X"BA",X"B6",X"BB",X"AB",X"62",X"48",X"47",
		X"44",X"48",X"42",X"7D",X"B3",X"B4",X"BA",X"B6",X"BB",X"AC",X"63",X"48",X"47",X"43",X"48",X"42",
		X"7C",X"B3",X"B4",X"BA",X"B6",X"BB",X"AD",X"64",X"48",X"47",X"43",X"48",X"41",X"79",X"B2",X"B4",
		X"BA",X"B6",X"BA",X"AF",X"66",X"47",X"48",X"43",X"48",X"40",X"77",X"B1",X"B5",X"BA",X"B7",X"BA",
		X"B1",X"69",X"47",X"48",X"42",X"48",X"40",X"74",X"B1",X"B5",X"BA",X"B8",X"BA",X"B3",X"6D",X"47",
		X"48",X"42",X"48",X"3F",X"6E",X"AF",X"B5",X"BA",X"B8",X"B9",X"B6",X"72",X"47",X"48",X"41",X"48",
		X"3F",X"68",X"AC",X"B6",X"B9",X"B9",X"B8",X"B8",X"79",X"47",X"48",X"41",X"48",X"3F",X"62",X"A9",
		X"B6",X"B9",X"B9",X"B7",X"BA",X"7F",X"49",X"49",X"42",X"48",X"40",X"5D",X"A5",X"B6",X"B8",X"BA",
		X"B6",X"BC",X"87",X"4B",X"49",X"42",X"48",X"41",X"56",X"A0",X"B7",X"B7",X"BA",X"B5",X"BC",X"8E",
		X"4D",X"49",X"42",X"47",X"43",X"50",X"99",X"B7",X"B6",X"BB",X"B5",X"BD",X"97",X"51",X"48",X"44",
		X"46",X"45",X"4A",X"91",X"B7",X"B6",X"BB",X"B6",X"BD",X"A1",X"58",X"47",X"45",X"44",X"46",X"45",
		X"86",X"B6",X"B5",X"BB",X"B5",X"BB",X"AA",X"61",X"47",X"47",X"43",X"48",X"42",X"79",X"B3",X"B5",
		X"BA",X"B6",X"B8",X"B1",X"6C",X"46",X"48",X"42",X"49",X"40",X"6C",X"AE",X"B6",X"B9",X"B8",X"B7",
		X"B7",X"78",X"47",X"49",X"42",X"49",X"41",X"60",X"A7",X"B6",X"B8",X"B9",X"B6",X"BB",X"86",X"4B",
		X"4A",X"43",X"49",X"43",X"55",X"9D",X"B6",X"B6",X"B9",X"B4",X"BC",X"94",X"50",X"49",X"44",X"47",
		X"45",X"4B",X"90",X"B6",X"B5",X"BA",X"B4",X"BC",X"A0",X"58",X"48",X"45",X"45",X"46",X"47",X"8A",
		X"B5",X"B5",X"BB",X"B5",X"BC",X"A2",X"5A",X"48",X"46",X"45",X"47",X"44",X"82",X"B4",X"B4",X"B9",
		X"B5",X"BA",X"AD",X"66",X"48",X"49",X"44",X"4A",X"41",X"72",X"B0",X"B5",X"B9",X"B7",X"B7",X"B6",
		X"74",X"47",X"49",X"42",X"49",X"40",X"61",X"A7",X"B5",X"B7",X"B9",X"B6",X"BC",X"87",X"4B",X"4A",
		X"43",X"48",X"42",X"52",X"9B",X"B6",X"B6",X"BA",X"B5",X"BD",X"99",X"54",X"49",X"45",X"46",X"46",
		X"47",X"8A",X"B5",X"B4",X"BA",X"B5",X"BB",X"A9",X"61",X"48",X"48",X"43",X"48",X"40",X"75",X"B0",
		X"B4",X"B9",X"B7",X"B8",X"B6",X"75",X"47",X"49",X"42",X"49",X"40",X"5F",X"A6",X"B6",X"B8",X"BA",
		X"B6",X"BD",X"8A",X"4C",X"49",X"43",X"47",X"42",X"4F",X"97",X"B6",X"B5",X"BB",X"B5",X"BD",X"9F",
		X"57",X"48",X"46",X"44",X"46",X"43",X"82",X"B4",X"B5",X"BA",X"B6",X"BB",X"B0",X"69",X"47",X"48",
		X"42",X"48",X"3F",X"6B",X"AD",X"B5",X"B9",X"B9",X"B8",X"BA",X"7D",X"49",X"49",X"42",X"48",X"40",
		X"58",X"A0",X"B7",X"B7",X"BB",X"B6",X"BD",X"95",X"51",X"49",X"44",X"45",X"45",X"48",X"8C",X"B6",
		X"B5",X"BB",X"B6",X"BC",X"AA",X"61",X"47",X"47",X"42",X"48",X"40",X"72",X"B0",X"B5",X"BA",X"B8",
		X"B8",X"B8",X"7A",X"48",X"49",X"41",X"48",X"41",X"59",X"A2",X"B7",X"B7",X"BB",X"B5",X"BD",X"95",
		X"51",X"48",X"44",X"45",X"45",X"47",X"8A",X"B6",X"B6",X"BB",X"B6",X"BB",X"AC",X"64",X"46",X"47",
		X"42",X"49",X"40",X"6D",X"AE",X"B6",X"B9",X"B8",X"B6",X"B9",X"80",X"48",X"48",X"42",X"48",X"42",
		X"52",X"9B",X"B8",X"B6",X"BB",X"B5",X"BD",X"9E",X"56",X"47",X"45",X"44",X"48",X"43",X"7F",X"B5",
		X"B6",X"BA",X"B7",X"B9",X"B3",X"70",X"46",X"49",X"42",X"49",X"40",X"60",X"A7",X"B7",X"B7",X"BA",
		X"B5",X"BC",X"90",X"4E",X"48",X"44",X"46",X"45",X"49",X"8C",X"B6",X"B5",X"BB",X"B5",X"BA",X"AC",
		X"64",X"46",X"48",X"43",X"4A",X"41",X"6B",X"AD",X"B6",X"B8",X"B9",X"B6",X"BA",X"85",X"4A",X"49",
		X"43",X"48",X"44",X"4E",X"95",X"B7",X"B5",X"BA",X"B4",X"BB",X"A5",X"5D",X"47",X"47",X"43",X"49",
		X"41",X"73",X"B0",X"B5",X"B9",X"B7",X"B6",X"B8",X"7D",X"49",X"4A",X"43",X"49",X"43",X"54",X"9B",
		X"B7",X"B5",X"BA",X"B4",X"BC",X"A0",X"58",X"48",X"47",X"44",X"48",X"42",X"7A",X"B2",X"B4",X"B9",
		X"B7",X"B7",X"B6",X"77",X"48",X"4A",X"42",X"49",X"41",X"57",X"9F",X"B6",X"B6",X"BA",X"B4",X"BD",
		X"9B",X"55",X"48",X"46",X"45",X"47",X"43",X"7E",X"B3",X"B4",X"B9",X"B7",X"B9",X"B6",X"74",X"48",
		X"4A",X"42",X"49",X"40",X"5A",X"A1",X"B6",X"B6",X"BA",X"B5",X"BD",X"9A",X"54",X"48",X"45",X"45",
		X"47",X"43",X"7E",X"B3",X"B4",X"BA",X"B7",X"B9",X"B6",X"74",X"48",X"49",X"42",X"49",X"40",X"58",
		X"A0",X"B6",X"B6",X"BA",X"B5",X"BD",X"9C",X"56",X"48",X"46",X"44",X"47",X"42",X"7B",X"B3",X"B5",
		X"BA",X"B8",X"B9",X"B8",X"79",X"48",X"4A",X"42",X"48",X"41",X"54",X"9D",X"B7",X"B6",X"BB",X"B5",
		X"BD",X"A1",X"59",X"47",X"46",X"43",X"47",X"40",X"74",X"B1",X"B5",X"B9",X"B8",X"B8",X"BA",X"80",
		X"49",X"49",X"42",X"47",X"42",X"4E",X"95",X"B7",X"B6",X"BB",X"B6",X"BD",X"A9",X"61",X"47",X"47",
		X"42",X"48",X"3F",X"6A",X"AC",X"B6",X"B9",X"BA",X"B6",X"BC",X"8C",X"4C",X"48",X"43",X"45",X"44",
		X"47",X"8A",X"B6",X"B5",X"BB",X"B7",X"BA",X"B1",X"6C",X"46",X"48",X"41",X"49",X"40",X"5D",X"A4",
		X"B7",X"B7",X"BB",X"B6",X"BD",X"9A",X"54",X"47",X"45",X"43",X"47",X"42",X"7B",X"B3",X"B6",X"BA",
		X"B8",X"B7",X"B8",X"7C",X"47",X"48",X"41",X"47",X"42",X"50",X"97",X"B7",X"B6",X"BB",X"B5",X"BC",
		X"A8",X"60",X"46",X"47",X"42",X"49",X"40",X"68",X"AC",X"B7",X"B8",X"BA",X"B6",X"BC",X"90",X"4E",
		X"48",X"44",X"45",X"46",X"46",X"85",X"B6",X"B5",X"BA",X"B6",X"B8",X"B4",X"73",X"46",X"49",X"42",
		X"49",X"41",X"56",X"9E",X"B8",X"B6",X"BB",X"B4",X"BC",X"A3",X"5B",X"46",X"47",X"43",X"49",X"41",
		X"6F",X"AF",X"B6",X"B8",X"B9",X"B5",X"BB",X"8A",X"4C",X"49",X"43",X"46",X"46",X"48",X"89",X"B6",
		X"B5",X"BA",X"B6",X"B8",X"B3",X"70",X"46",X"49",X"42",X"49",X"42",X"57",X"9F",X"B7",X"B6",X"BA",
		X"B4",X"BC",X"A2",X"5B",X"47",X"47",X"43",X"4A",X"41",X"6D",X"AE",X"B6",X"B8",X"B9",X"B5",X"BC",
		X"8D",X"4D",X"49",X"44",X"46",X"47",X"46",X"85",X"B5",X"B5",X"BA",X"B6",X"B8",X"B5",X"76",X"47",
		X"4A",X"43",X"49",X"42",X"52",X"9A",X"B7",X"B5",X"BA",X"B4",X"BB",X"A9",X"62",X"46",X"48",X"43",
		X"4A",X"40",X"64",X"A8",X"B6",X"B6",X"B9",X"B5",X"BD",X"97",X"53",X"48",X"46",X"45",X"48",X"42",
		X"78",X"B1",X"B5",X"B8",X"B8",X"B7",X"BB",X"85",X"4B",X"4A",X"44",X"47",X"45",X"49",X"8C",X"B6",
		X"B4",X"BA",X"B6",X"B9",X"B2",X"6F",X"47",X"4A",X"42",X"49",X"41",X"56",X"9D",X"B6",X"B5",X"BA",
		X"B5",X"BC",X"A6",X"5E",X"47",X"48",X"42",X"49",X"3F",X"67",X"AA",X"B6",X"B7",X"BA",X"B6",X"BD",
		X"96",X"53",X"48",X"45",X"44",X"47",X"41",X"78",X"B1",X"B5",X"B9",X"B8",X"B7",X"BC",X"87",X"4B",
		X"49",X"44",X"46",X"45",X"46",X"87",X"B5",X"B5",X"BA",X"B7",X"B9",X"B6",X"76",X"47",X"49",X"42",
		X"48",X"42",X"50",X"96",X"B7",X"B6",X"BB",X"B6",X"BB",X"AC",X"64",X"45",X"47",X"41",X"48",X"3F",
		X"62",X"A8",X"B7",X"B8",X"BB",X"B6",X"BE",X"95",X"52",X"48",X"45",X"44",X"46",X"41",X"7A",X"B2",
		X"B5",X"B9",X"B9",X"B7",X"BB",X"85",X"4B",X"49",X"43",X"46",X"44",X"46",X"88",X"B6",X"B5",X"BB",
		X"B7",X"B9",X"B6",X"77",X"47",X"49",X"42",X"47",X"42",X"4E",X"94",X"B8",X"B6",X"BC",X"B6",X"BB",
		X"B0",X"6A",X"45",X"48",X"41",X"48",X"40",X"57",X"9F",X"B8",X"B7",X"BC",X"B6",X"BD",X"A7",X"5F",
		X"46",X"47",X"41",X"49",X"3F",X"62",X"A8",X"B7",X"B7",X"BB",X"B5",X"BD",X"9E",X"57",X"46",X"46",
		X"42",X"48",X"40",X"6C",X"AD",X"B7",X"B9",X"BA",X"B5",X"BD",X"95",X"51",X"47",X"45",X"43",X"48",
		X"41",X"75",X"B1",X"B7",X"B9",X"B9",X"B6",X"BC",X"8E",X"4D",X"47",X"44",X"44",X"47",X"43",X"7C",
		X"B4",X"B6",X"BA",X"B9",X"B7",X"BB",X"87",X"4B",X"48",X"43",X"45",X"46",X"45",X"83",X"B5",X"B6",
		X"BA",X"B8",X"B7",X"B9",X"7F",X"48",X"48",X"43",X"47",X"45",X"48",X"8A",X"B7",X"B5",X"BA",X"B7",
		X"B8",X"B6",X"78",X"47",X"49",X"42",X"48",X"44",X"4C",X"90",X"B7",X"B5",X"BA",X"B6",X"B9",X"B3",
		X"73",X"46",X"49",X"42",X"48",X"43",X"4F",X"95",X"B8",X"B5",X"BB",X"B6",X"B9",X"B1",X"6E",X"46",
		X"49",X"41",X"49",X"42",X"51",X"98",X"B7",X"B5",X"BB",X"B5",X"BA",X"B0",X"6C",X"46",X"49",X"42",
		X"49",X"42",X"52",X"99",X"B8",X"B5",X"BA",X"B5",X"BA",X"AF",X"6B",X"46",X"49",X"42",X"49",X"42",
		X"53",X"9A",X"B7",X"B5",X"BA",X"B5",X"BA",X"AF",X"6B",X"46",X"49",X"42",X"4A",X"42",X"54",X"9A",
		X"B7",X"B5",X"BA",X"B5",X"BB",X"AF",X"6A",X"46",X"49",X"42",X"49",X"42",X"54",X"9B",X"B7",X"B5",
		X"BA",X"B5",X"BB",X"AE",X"6A",X"46",X"49",X"42",X"49",X"41",X"54",X"9B",X"B7",X"B5",X"BA",X"B5",
		X"BB",X"AF",X"6A",X"46",X"49",X"42",X"49",X"41",X"53",X"99",X"B7",X"B5",X"BB",X"B5",X"BB",X"B0",
		X"6C",X"46",X"4A",X"42",X"49",X"41",X"52",X"98",X"B7",X"B5",X"BB",X"B6",X"BB",X"B1",X"6E",X"46",
		X"49",X"42",X"49",X"42",X"50",X"96",X"B7",X"B5",X"BB",X"B6",X"BB",X"B3",X"70",X"47",X"4A",X"42",
		X"48",X"42",X"4E",X"93",X"B7",X"B5",X"BB",X"B6",X"BA",X"B4",X"73",X"47",X"4A",X"42",X"48",X"43",
		X"4B",X"90",X"B7",X"B5",X"BB",X"B7",X"B9",X"B6",X"78",X"47",X"49",X"42",X"47",X"43",X"48",X"8B",
		X"B6",X"B5",X"BA",X"B7",X"B9",X"B9",X"7E",X"48",X"49",X"43",X"46",X"44",X"45",X"85",X"B5",X"B5",
		X"BA",X"B8",X"B8",X"BB",X"85",X"4A",X"48",X"43",X"45",X"46",X"43",X"7D",X"B3",X"B6",X"BA",X"B9",
		X"B7",X"BD",X"8D",X"4E",X"48",X"44",X"44",X"47",X"41",X"75",X"B1",X"B6",X"B9",X"BA",X"B6",X"BD",
		X"95",X"52",X"47",X"45",X"42",X"48",X"3F",X"6C",X"AD",X"B7",X"B8",X"BB",X"B6",X"BD",X"9D",X"57",
		X"46",X"46",X"41",X"48",X"3F",X"63",X"A8",X"B7",X"B7",X"BB",X"B5",X"BD",X"A5",X"5E",X"45",X"47",
		X"41",X"49",X"40",X"5B",X"A1",X"B8",X"B6",X"BC",X"B5",X"BC",X"AD",X"67",X"45",X"48",X"41",X"49",
		X"41",X"52",X"99",X"B8",X"B6",X"BC",X"B6",X"BA",X"B4",X"72",X"46",X"48",X"41",X"47",X"43",X"4B",
		X"8E",X"B8",X"B6",X"BB",X"B7",X"B8",X"B8",X"7F",X"48",X"48",X"43",X"46",X"46",X"45",X"81",X"B5",
		X"B6",X"BA",X"B9",X"B6",X"BC",X"8C",X"4D",X"47",X"44",X"44",X"48",X"40",X"72",X"B0",X"B7",X"B8",
		X"BA",X"B5",X"BC",X"9A",X"55",X"46",X"47",X"42",X"49",X"40",X"63",X"A7",X"B8",X"B7",X"BB",X"B5",
		X"BC",X"A8",X"61",X"45",X"48",X"42",X"4A",X"42",X"55",X"9C",X"B8",X"B6",X"BB",X"B6",X"BA",X"B3",
		X"71",X"46",X"49",X"42",X"48",X"44",X"4A",X"8C",X"B7",X"B5",X"BA",X"B7",X"B6",X"B9",X"83",X"4A",
		X"48",X"44",X"45",X"47",X"43",X"7A",X"B3",X"B6",X"B8",X"B8",X"B4",X"BC",X"95",X"52",X"46",X"46",
		X"43",X"49",X"40",X"66",X"A9",X"B7",X"B6",X"BA",X"B4",X"BC",X"A6",X"60",X"45",X"49",X"42",X"4A",
		X"41",X"55",X"9B",X"B8",X"B5",X"BA",X"B5",X"B9",X"B3",X"73",X"46",X"4A",X"43",X"48",X"45",X"49",
		X"89",X"B6",X"B5",X"B9",X"B8",X"B7",X"BB",X"88",X"4C",X"49",X"45",X"45",X"48",X"41",X"73",X"B0",
		X"B6",X"B7",X"B9",X"B4",X"BD",X"9D",X"58",X"47",X"48",X"43",X"4A",X"40",X"5E",X"A3",X"B7",X"B5",
		X"BA",X"B5",X"BB",X"AE",X"69",X"46",X"4A",X"42",X"48",X"42",X"4D",X"91",X"B6",X"B4",X"BA",X"B7",
		X"B8",X"B9",X"80",X"4A",X"49",X"44",X"46",X"47",X"42",X"7A",X"B2",X"B5",X"B8",X"B9",X"B6",X"BD",
		X"98",X"54",X"47",X"47",X"43",X"49",X"3F",X"62",X"A6",X"B7",X"B6",X"BB",X"B5",X"BC",X"AC",X"66",
		X"46",X"49",X"41",X"48",X"41",X"4E",X"93",X"B7",X"B5",X"BA",X"B7",X"B9",X"B9",X"7E",X"49",X"49",
		X"43",X"45",X"46",X"42",X"7A",X"B2",X"B6",X"B8",X"BA",X"B6",X"BE",X"98",X"54",X"47",X"47",X"42",
		X"49",X"3F",X"60",X"A5",X"B7",X"B6",X"BB",X"B6",X"BC",X"AE",X"69",X"45",X"49",X"41",X"48",X"42",
		X"4B",X"8F",X"B7",X"B6",X"BB",X"B8",X"B8",X"BB",X"85",X"4B",X"48",X"44",X"44",X"47",X"40",X"73",
		X"B0",X"B7",X"B8",X"BA",X"B5",X"BD",X"A0",X"59",X"45",X"47",X"41",X"48",X"3F",X"58",X"9F",X"B8",
		X"B6",X"BB",X"B6",X"BA",X"B4",X"73",X"46",X"48",X"42",X"46",X"45",X"45",X"84",X"B5",X"B6",X"BA",
		X"BA",X"B6",X"BD",X"92",X"50",X"46",X"45",X"42",X"49",X"40",X"64",X"A9",X"B8",X"B8",X"BC",X"B6",
		X"BC",X"AD",X"67",X"45",X"48",X"41",X"47",X"43",X"4B",X"8F",X"B8",X"B7",X"BB",X"B8",X"B7",X"BB",
		X"88",X"4B",X"47",X"44",X"43",X"48",X"40",X"6D",X"AE",X"B8",X"B8",X"BB",X"B5",X"BC",X"A7",X"60",
		X"45",X"47",X"41",X"48",X"42",X"50",X"96",X"B8",X"B6",X"BB",X"B7",X"B7",X"B9",X"80",X"49",X"47",
		X"44",X"45",X"48",X"42",X"74",X"B1",X"B7",X"B8",X"BA",X"B5",X"BC",X"A2",X"5B",X"45",X"47",X"42",
		X"49",X"42",X"54",X"9B",X"B8",X"B6",X"BA",X"B7",X"B8",X"B8",X"7C",X"48",X"48",X"44",X"45",X"48",
		X"43",X"78",X"B2",X"B7",X"B8",X"B9",X"B4",X"BC",X"9F",X"59",X"46",X"47",X"42",X"49",X"42",X"55",
		X"9C",X"B8",X"B6",X"BA",X"B6",X"B7",X"B7",X"7B",X"48",X"48",X"44",X"46",X"48",X"42",X"78",X"B2",
		X"B6",X"B8",X"B9",X"B5",X"BC",X"A1",X"5A",X"46",X"47",X"43",X"49",X"42",X"54",X"9B",X"B7",X"B6",
		X"BA",X"B7",X"B7",X"B9",X"7D",X"49",X"48",X"44",X"45",X"47",X"41",X"75",X"B0",X"B6",X"B7",X"B9",
		X"B5",X"BC",X"A3",X"5C",X"46",X"48",X"43",X"49",X"42",X"51",X"98",X"B7",X"B6",X"B9",X"B7",X"B7",
		X"B9",X"80",X"4A",X"48",X"45",X"45",X"48",X"41",X"71",X"AF",X"B6",X"B7",X"B9",X"B5",X"BB",X"A7",
		X"60",X"47",X"48",X"44",X"48",X"44",X"4C",X"92",X"B6",X"B6",X"B9",X"B8",X"B6",X"BC",X"8B",X"4E",
		X"48",X"46",X"44",X"49",X"41",X"65",X"AA",X"B6",X"B7",X"B9",X"B6",X"B9",X"B0",X"6A",X"47",X"48",
		X"44",X"46",X"46",X"45",X"85",X"B4",X"B6",X"B8",X"B9",X"B6",X"BC",X"99",X"54",X"48",X"46",X"44",
		X"48",X"42",X"56",X"9F",X"B5",X"B7",X"B9",X"B8",X"B8",X"BA",X"7D",X"4A",X"48",X"45",X"45",X"48",
		X"41",X"70",X"AF",X"B5",X"B8",X"B9",X"B7",X"BB",X"AC",X"63",X"48",X"47",X"44",X"46",X"45",X"49",
		X"8D",X"B5",X"B6",X"B9",X"B8",X"B6",X"BC",X"91",X"50",X"48",X"45",X"44",X"47",X"40",X"5D",X"A5",
		X"B6",X"B7",X"B9",X"B7",X"B8",X"B6",X"74",X"48",X"48",X"43",X"45",X"46",X"42",X"79",X"B2",X"B6",
		X"B9",X"BA",X"B7",X"BE",X"9D",X"56",X"46",X"46",X"42",X"47",X"40",X"59",X"A2",X"B6",X"B8",X"BA",
		X"B9",X"B9",X"B9",X"7A",X"4A",X"48",X"44",X"44",X"47",X"40",X"70",X"AF",X"B5",X"B8",X"B9",X"B7",
		X"BA",X"AB",X"61",X"47",X"46",X"43",X"45",X"45",X"47",X"8C",X"B5",X"B7",X"B9",X"BA",X"B6",X"BC",
		X"94",X"50",X"47",X"44",X"44",X"47",X"42",X"58",X"A3",X"B6",X"B9",X"B9",X"BA",X"B7",X"BA",X"7C",
		X"49",X"46",X"44",X"44",X"47",X"41",X"6E",X"B0",X"B6",X"BA",X"B9",X"B9",X"B9",X"B0",X"66",X"48",
		X"45",X"44",X"44",X"46",X"44",X"84",X"B5",X"B7",X"BA",X"B9",X"B6",X"BB",X"9F",X"56",X"47",X"44",
		X"44",X"45",X"44",X"4D",X"98",X"B6",X"B8",X"B9",X"BA",X"B5",X"BC",X"8B",X"4C",X"47",X"44",X"44",
		X"47",X"42",X"5E",X"A8",X"B6",X"BA",X"B8",X"BA",X"B6",X"B8",X"75",X"49",X"46",X"44",X"44",X"48",
		X"42",X"71",X"B1",X"B6",X"BA",X"B8",X"B8",X"B8",X"AE",X"63",X"48",X"45",X"45",X"44",X"47",X"45",
		X"86",X"B5",X"B7",X"B9",X"B8",X"B6",X"BA",X"A0",X"55",X"48",X"44",X"45",X"45",X"46",X"4C",X"97",
		X"B5",X"B8",X"B8",X"B9",X"B5",X"BB",X"90",X"4E",X"48",X"44",X"45",X"47",X"44",X"57",X"A4",X"B5",
		X"BA",X"B7",X"BA",X"B5",X"BA",X"7E",X"4A",X"47",X"45",X"45",X"48",X"43",X"66",X"AD",X"B5",X"BA",
		X"B7",X"B9",X"B6",X"B6",X"6F",X"49",X"46",X"45",X"44",X"48",X"42",X"76",X"B2",X"B5",X"BA",X"B7",
		X"B7",X"B7",X"AD",X"60",X"48",X"45",X"46",X"44",X"48",X"44",X"86",X"B4",X"B6",X"B9",X"B8",X"B6",
		X"BA",X"A2",X"57",X"49",X"44",X"46",X"45",X"47",X"4A",X"93",X"B5",X"B8",X"B8",X"B9",X"B5",X"BC",
		X"97",X"51",X"49",X"44",X"47",X"46",X"46",X"50",X"9E",X"B4",X"B9",X"B7",X"B9",X"B5",X"BC",X"8B",
		X"4D",X"49",X"45",X"46",X"47",X"44",X"58",X"A5",X"B4",X"B9",X"B6",X"B9",X"B4",X"BB",X"80",X"4B",
		X"48",X"45",X"45",X"47",X"42",X"61",X"AA",X"B3",X"BA",X"B6",X"BA",X"B5",X"B9",X"76",X"4A",X"47",
		X"46",X"45",X"48",X"42",X"69",X"AE",X"B3",X"BA",X"B6",X"BA",X"B6",X"B7",X"6E",X"4A",X"46",X"46",
		X"44",X"48",X"41",X"72",X"B1",X"B4",X"BA",X"B7",X"B9",X"B7",X"B3",X"67",X"4A",X"46",X"46",X"44",
		X"48",X"42",X"79",X"B2",X"B5",X"BA",X"B7",X"B8",X"B8",X"AF",X"62",X"4A",X"45",X"46",X"43",X"47",
		X"42",X"80",X"B3",X"B5",X"B9",X"B8",X"B8",X"B9",X"AB",X"5D",X"4A",X"44",X"46",X"43",X"47",X"43",
		X"86",X"B3",X"B6",X"B9",X"B8",X"B8",X"BA",X"A6",X"59",X"4A",X"44",X"46",X"44",X"47",X"45",X"8B",
		X"B4",X"B7",X"B9",X"B9",X"B7",X"BB",X"A3",X"57",X"49",X"44",X"46",X"44",X"47",X"46",X"8F",X"B4",
		X"B7",X"B9",X"B9",X"B7",X"BC",X"A0",X"55",X"49",X"43",X"45",X"43",X"46",X"48",X"92",X"B4",X"B8",
		X"B8",X"BA",X"B7",X"BC",X"9D",X"53",X"49",X"43",X"45",X"43",X"45",X"49",X"94",X"B4",X"B8",X"B8",
		X"BA",X"B6",X"BC",X"9B",X"52",X"49",X"43",X"46",X"43",X"46",X"49",X"95",X"B4",X"B9",X"B9",X"BA",
		X"B7",X"BC",X"9B",X"52",X"49",X"43",X"46",X"44",X"46",X"4A",X"96",X"B5",X"B9",X"B9",X"BB",X"B7",
		X"BD",X"9B",X"53",X"49",X"43",X"46",X"44",X"46",X"49",X"95",X"B5",X"B9",X"B9",X"BA",X"B7",X"BC",
		X"9D",X"53",X"49",X"43",X"45",X"43",X"47",X"49",X"93",X"B5",X"B8",X"B9",X"B9",X"B6",X"BB",X"9F",
		X"54",X"48",X"42",X"45",X"43",X"47",X"46",X"8E",X"B5",X"B8",X"B9",X"B9",X"B7",X"BA",X"A4",X"57",
		X"48",X"43",X"46",X"43",X"48",X"45",X"89",X"B5",X"B7",X"BA",X"B8",X"B7",X"B9",X"A8",X"5A",X"48",
		X"43",X"46",X"44",X"48",X"44",X"84",X"B5",X"B7",X"BA",X"B8",X"B8",X"B8",X"AD",X"5F",X"48",X"43",
		X"46",X"43",X"48",X"43",X"7C",X"B4",X"B6",X"BB",X"B7",X"B9",X"B7",X"B1",X"65",X"49",X"44",X"46",
		X"44",X"48",X"42",X"75",X"B3",X"B5",X"BB",X"B6",X"B9",X"B6",X"B5",X"6B",X"49",X"45",X"45",X"44",
		X"48",X"42",X"6D",X"B0",X"B4",X"BB",X"B6",X"BA",X"B4",X"B8",X"73",X"49",X"46",X"44",X"44",X"47",
		X"42",X"63",X"AC",X"B4",X"BB",X"B6",X"BA",X"B3",X"BA",X"7D",X"4A",X"47",X"44",X"45",X"47",X"44",
		X"5A",X"A7",X"B4",X"BA",X"B6",X"BA",X"B4",X"BC",X"88",X"4C",X"48",X"44",X"46",X"46",X"46",X"52",
		X"9F",X"B4",X"B9",X"B7",X"BA",X"B5",X"BC",X"94",X"50",X"49",X"44",X"47",X"45",X"47",X"4B",X"96",
		X"B5",X"B8",X"B8",X"B9",X"B6",X"BB",X"A0",X"56",X"49",X"44",X"47",X"45",X"48",X"45",X"8A",X"B5",
		X"B6",X"B9",X"B7",X"B7",X"B9",X"AB",X"5E",X"4A",X"45",X"47",X"44",X"49",X"42",X"7A",X"B3",X"B5",
		X"BA",X"B6",X"B9",X"B6",X"B5",X"6A",X"4A",X"46",X"46",X"44",X"48",X"41",X"69",X"AF",X"B3",X"BA",
		X"B5",X"BA",X"B4",X"BA",X"7A",X"4B",X"48",X"45",X"45",X"46",X"43",X"59",X"A6",X"B3",X"B9",X"B6",
		X"BA",X"B4",X"BC",X"8D",X"4E",X"49",X"44",X"46",X"45",X"46",X"4C",X"99",X"B4",X"B8",X"B8",X"B9",
		X"B6",X"BB",X"9F",X"55",X"4A",X"44",X"47",X"44",X"47",X"44",X"87",X"B4",X"B6",X"B9",X"B8",X"B9",
		X"B9",X"AF",X"62",X"4A",X"45",X"46",X"44",X"48",X"41",X"72",X"B1",X"B4",X"BB",X"B6",X"BA",X"B6",
		X"BA",X"75",X"4A",X"47",X"45",X"44",X"47",X"42",X"5D",X"A9",X"B3",X"BA",X"B6",X"BB",X"B5",X"BE",
		X"8B",X"4D",X"48",X"43",X"45",X"44",X"45",X"4C",X"99",X"B4",X"B8",X"B8",X"B9",X"B6",X"BC",X"A1",
		X"56",X"49",X"43",X"46",X"43",X"47",X"43",X"84",X"B4",X"B6",X"BA",X"B8",X"B9",X"B8",X"B2",X"66",
		X"49",X"45",X"45",X"43",X"47",X"41",X"6B",X"AF",X"B4",X"BB",X"B7",X"BB",X"B5",X"BB",X"7C",X"4A",
		X"47",X"44",X"45",X"45",X"43",X"55",X"A3",X"B4",X"BA",X"B8",X"BB",X"B6",X"BD",X"96",X"50",X"49",
		X"43",X"46",X"43",X"46",X"47",X"8E",X"B5",X"B7",X"BA",X"B9",X"B9",X"B9",X"AC",X"5E",X"49",X"44",
		X"45",X"43",X"48",X"41",X"73",X"B2",X"B5",X"BC",X"B7",X"BB",X"B6",X"BA",X"77",X"49",X"46",X"44",
		X"44",X"46",X"43",X"59",X"A6",X"B5",X"BB",X"B8",X"BB",X"B5",X"BD",X"94",X"4F",X"48",X"42",X"45",
		X"44",X"47",X"47",X"8F",X"B5",X"B8",X"BA",X"B9",X"B8",X"B9",X"AD",X"60",X"48",X"44",X"45",X"43",
		X"48",X"42",X"70",X"B2",X"B5",X"BC",X"B7",X"BB",X"B5",X"BB",X"7B",X"49",X"46",X"43",X"45",X"45",
		X"44",X"54",X"A2",X"B5",X"BA",X"B8",X"BA",X"B5",X"BB",X"9A",X"52",X"48",X"43",X"46",X"43",X"48",
		X"44",X"86",X"B5",X"B6",X"BA",X"B7",X"B9",X"B7",X"B2",X"67",X"48",X"45",X"45",X"44",X"48",X"42",
		X"66",X"AE",X"B5",X"BB",X"B7",X"BB",X"B4",X"BC",X"86",X"4A",X"47",X"42",X"45",X"44",X"46",X"4C",
		X"98",X"B5",X"B8",X"B9",X"B9",X"B7",X"BA",X"A7",X"5A",X"48",X"43",X"46",X"44",X"49",X"42",X"77",
		X"B3",X"B5",X"BB",X"B7",X"BA",X"B5",X"B9",X"76",X"49",X"47",X"44",X"45",X"47",X"45",X"57",X"A4",
		X"B5",X"BA",X"B7",X"B9",X"B5",X"BB",X"9B",X"53",X"49",X"44",X"47",X"44",X"49",X"44",X"82",X"B5",
		X"B6",X"BA",X"B6",X"B8",X"B5",X"B5",X"6D",X"49",X"46",X"45",X"45",X"48",X"43",X"5D",X"A9",X"B4",
		X"BA",X"B6",X"BA",X"B4",X"BC",X"92",X"4F",X"49",X"44",X"47",X"45",X"48",X"46",X"89",X"B5",X"B6",
		X"B9",X"B7",X"B8",X"B6",X"B3",X"68",X"49",X"46",X"46",X"45",X"48",X"43",X"61",X"AB",X"B4",X"BA",
		X"B6",X"BA",X"B4",X"BC",X"8F",X"4E",X"49",X"44",X"47",X"45",X"48",X"47",X"8C",X"B5",X"B6",X"BA",
		X"B7",X"B8",X"B7",X"B2",X"68",X"49",X"46",X"46",X"45",X"48",X"42",X"61",X"AB",X"B3",X"BA",X"B6",
		X"BA",X"B4",X"BD",X"91",X"4F",X"49",X"44",X"47",X"44",X"47",X"46",X"8B",X"B4",X"B5",X"B9",X"B7",
		X"B8",X"B7",X"B2",X"68",X"4A",X"46",X"46",X"45",X"47",X"42",X"61",X"AB",X"B3",X"B9",X"B5",X"BA",
		X"B4",X"BC",X"91",X"4F",X"49",X"44",X"47",X"45",X"48",X"46",X"89",X"B4",X"B5",X"B9",X"B6",X"B8",
		X"B6",X"B3",X"6A",X"48",X"46",X"45",X"45",X"46",X"43",X"5B",X"A7",X"B3",X"BA",X"B6",X"BB",X"B5",
		X"BD",X"97",X"53",X"48",X"44",X"45",X"45",X"45",X"4B",X"95",X"B5",X"B8",X"B9",X"BA",X"B7",X"BD",
		X"9A",X"53",X"4A",X"43",X"47",X"43",X"48",X"42",X"80",X"B3",X"B5",X"BA",X"B7",X"BA",X"B6",X"B9",
		X"75",X"4B",X"47",X"45",X"45",X"46",X"43",X"52",X"9F",X"B4",X"B8",X"B7",X"B9",X"B6",X"BB",X"A5",
		X"5A",X"4A",X"44",X"46",X"44",X"48",X"41",X"70",X"B0",X"B4",X"BB",X"B6",X"BB",X"B4",X"BC",X"84",
		X"4C",X"48",X"44",X"46",X"44",X"46",X"48",X"92",X"B5",X"B7",X"BA",X"B9",X"B9",X"B8",X"B1",X"65",
		X"49",X"45",X"45",X"44",X"47",X"41",X"60",X"AA",X"B4",X"BB",X"B7",X"BB",X"B6",X"BE",X"97",X"51",
		X"49",X"43",X"46",X"43",X"47",X"42",X"7E",X"B4",X"B5",X"BB",X"B7",X"BB",X"B6",X"BB",X"7B",X"4A",
		X"47",X"44",X"45",X"44",X"45",X"4D",X"98",X"B5",X"B8",X"B9",X"B9",X"B8",X"B9",X"AE",X"61",X"48",
		X"44",X"45",X"43",X"47",X"41",X"62",X"AB",X"B4",X"BB",X"B7",X"BB",X"B5",X"BD",X"96",X"50",X"48",
		X"42",X"45",X"43",X"47",X"42",X"7E",X"B4",X"B6",X"BC",X"B7",X"BB",X"B5",X"BA",X"7A",X"49",X"46",
		X"43",X"45",X"45",X"44",X"4F",X"9C",X"B5",X"B9",X"B9",X"BA",X"B7",X"BB",X"A6",X"59",X"48",X"43",
		X"45",X"43",X"48",X"41",X"6B",X"B0",X"B5",X"BC",X"B7",X"BB",X"B5",X"BD",X"90",X"4E",X"48",X"43",
		X"46",X"44",X"48",X"44",X"83",X"B5",X"B6",X"BB",X"B7",X"BA",X"B5",X"B9",X"78",X"49",X"46",X"43",
		X"45",X"45",X"45",X"4D",X"99",X"B6",X"B9",X"BA",X"B8",X"B8",X"B8",X"AF",X"63",X"48",X"44",X"45",
		X"44",X"47",X"43",X"5D",X"A9",X"B5",X"BB",X"B8",X"BA",X"B5",X"BB",X"9E",X"54",X"48",X"43",X"46",
		X"44",X"49",X"42",X"72",X"B2",X"B5",X"BC",X"B7",X"BB",X"B4",X"BC",X"8A",X"4C",X"48",X"43",X"46",
		X"44",X"48",X"45",X"85",X"B6",X"B6",X"BB",X"B7",X"BA",X"B5",X"B9",X"78",X"49",X"47",X"43",X"46",
		X"45",X"46",X"4C",X"96",X"B6",X"B8",X"B9",X"B7",X"B8",X"B7",X"B2",X"68",X"48",X"46",X"45",X"45",
		X"47",X"44",X"58",X"A4",X"B5",X"B9",X"B8",X"B9",X"B5",X"B9",X"A6",X"5A",X"48",X"44",X"46",X"44",
		X"48",X"42",X"66",X"AD",X"B4",X"BB",X"B6",X"BA",X"B4",X"BB",X"98",X"51",X"48",X"43",X"47",X"44",
		X"49",X"42",X"76",X"B3",X"B5",X"BB",X"B6",X"BA",X"B4",X"BC",X"89",X"4C",X"48",X"43",X"47",X"45",
		X"48",X"45",X"85",X"B5",X"B6",X"BB",X"B6",X"BA",X"B5",X"BA",X"78",X"49",X"47",X"44",X"46",X"45",
		X"46",X"4C",X"96",X"B5",X"B7",X"B9",X"B7",X"B7",X"B7",X"B2",X"68",X"49",X"46",X"45",X"45",X"47",
		X"43",X"55",X"A2",X"B4",X"B8",X"B7",X"B8",X"B6",X"B9",X"AA",X"5E",X"49",X"45",X"46",X"45",X"48",
		X"42",X"5E",X"A8",X"B4",X"B9",X"B6",X"B9",X"B5",X"BB",X"A2",X"58",X"49",X"45",X"47",X"45",X"49",
		X"42",X"67",X"AD",X"B4",X"BA",X"B6",X"BA",X"B5",X"BC",X"9B",X"53",X"49",X"44",X"47",X"44",X"49",
		X"42",X"70",X"B1",X"B4",X"BB",X"B6",X"BB",X"B4",X"BD",X"91",X"4F",X"49",X"44",X"47",X"44",X"48",
		X"42",X"79",X"B3",X"B4",X"BB",X"B6",X"BA",X"B4",X"BD",X"8A",X"4D",X"49",X"44",X"47",X"44",X"48",
		X"42",X"7E",X"B3",X"B4",X"BA",X"B6",X"BA",X"B4",X"BC",X"85",X"4C",X"49",X"44",X"47",X"44",X"47",
		X"44",X"84",X"B4",X"B4",X"BA",X"B6",X"BA",X"B5",X"BB",X"7E",X"4B",X"48",X"44",X"46",X"44",X"47",
		X"46",X"8A",X"B5",X"B6",X"BA",X"B7",X"BA",X"B6",X"BB",X"7A",X"4A",X"48",X"44",X"46",X"44",X"46",
		X"48",X"8F",X"B5",X"B6",X"BA",X"B7",X"BA",X"B7",X"BA",X"76",X"4A",X"47",X"44",X"45",X"44",X"45",
		X"48",X"91",X"B5",X"B6",X"BA",X"B7",X"BA",X"B7",X"B9",X"74",X"4A",X"47",X"44",X"46",X"44",X"45",
		X"49",X"93",X"B5",X"B6",X"B9",X"B7",X"B9",X"B6",X"B7",X"72",X"49",X"47",X"44",X"45",X"44",X"45",
		X"4A",X"93",X"B5",X"B7",X"BA",X"B7",X"B9",X"B6",X"B7",X"72",X"48",X"46",X"43",X"45",X"45",X"46",
		X"4A",X"93",X"B6",X"B7",X"BB",X"B8",X"BA",X"B6",X"B8",X"74",X"48",X"46",X"43",X"45",X"44",X"46",
		X"4A",X"91",X"B6",X"B8",X"BB",X"B8",X"BB",X"B7",X"B9",X"74",X"48",X"46",X"43",X"44",X"44",X"45",
		X"4D",X"98",X"B6",X"B9",X"BB",X"BA",X"BA",X"B9",X"B3",X"69",X"49",X"45",X"44",X"44",X"45",X"43",
		X"51",X"9E",X"B6",X"B8",X"BA",X"B9",X"B9",X"B8",X"B3",X"6A",X"49",X"46",X"44",X"44",X"45",X"44",
		X"4E",X"99",X"B6",X"B8",X"BA",X"B8",X"B9",X"B7",X"B6",X"6F",X"48",X"46",X"43",X"45",X"45",X"45",
		X"4A",X"93",X"B6",X"B7",X"BA",X"B7",X"B9",X"B5",X"B8",X"75",X"48",X"46",X"43",X"46",X"45",X"47",
		X"47",X"8D",X"B6",X"B7",X"BB",X"B7",X"BA",X"B5",X"BA",X"7C",X"49",X"47",X"43",X"46",X"44",X"48",
		X"46",X"87",X"B6",X"B6",X"BC",X"B7",X"BB",X"B4",X"BB",X"84",X"4A",X"47",X"42",X"46",X"44",X"48",
		X"43",X"7E",X"B5",X"B6",X"BC",X"B7",X"BB",X"B4",X"BC",X"8D",X"4D",X"48",X"43",X"46",X"43",X"49",
		X"42",X"75",X"B3",X"B5",X"BC",X"B6",X"BA",X"B4",X"BC",X"95",X"50",X"48",X"43",X"46",X"43",X"49",
		X"42",X"6C",X"B0",X"B5",X"BB",X"B6",X"BA",X"B4",X"BB",X"9F",X"56",X"48",X"44",X"46",X"44",X"48",
		X"42",X"61",X"AA",X"B5",X"BA",X"B7",X"B9",X"B5",X"B9",X"A9",X"5E",X"48",X"45",X"45",X"44",X"47",
		X"44",X"56",X"A2",X"B6",X"B9",X"B8",X"B8",X"B7",X"B7",X"B1",X"68",X"48",X"46",X"45",X"46",X"47",
		X"46",X"4D",X"97",X"B6",X"B7",X"B9",X"B6",X"B8",X"B4",X"B8",X"77",X"49",X"48",X"44",X"47",X"46",
		X"48",X"46",X"86",X"B5",X"B5",X"BA",X"B5",X"BA",X"B3",X"BC",X"89",X"4C",X"48",X"44",X"47",X"45",
		X"49",X"43",X"74",X"B2",X"B4",X"BB",X"B6",X"BA",X"B4",X"BC",X"9A",X"53",X"48",X"44",X"47",X"45",
		X"49",X"42",X"64",X"AC",X"B5",X"BA",X"B7",X"B9",X"B6",X"BA",X"A9",X"5D",X"48",X"45",X"46",X"45",
		X"47",X"44",X"56",X"A1",X"B5",X"B8",X"B8",X"B8",X"B8",X"B8",X"B4",X"6C",X"49",X"47",X"45",X"46",
		X"46",X"46",X"4A",X"92",X"B6",X"B6",X"BA",X"B6",X"BA",X"B5",X"BB",X"7E",X"4B",X"49",X"44",X"47",
		X"44",X"48",X"43",X"7E",X"B4",X"B4",X"BA",X"B5",X"BA",X"B4",X"BD",X"93",X"50",X"49",X"44",X"46",
		X"43",X"48",X"41",X"68",X"AD",X"B4",X"BA",X"B7",X"BA",X"B6",X"BB",X"A6",X"5B",X"48",X"44",X"45",
		X"43",X"46",X"42",X"57",X"A3",X"B4",X"B8",X"B8",X"B9",X"B8",X"B8",X"B2",X"69",X"49",X"46",X"44",
		X"45",X"45",X"44",X"4A",X"92",X"B5",X"B6",X"BA",X"B7",X"BA",X"B5",X"BB",X"80",X"4B",X"48",X"43",
		X"46",X"43",X"47",X"41",X"79",X"B3",X"B4",X"BB",X"B6",X"BB",X"B5",X"BD",X"99",X"53",X"49",X"44",
		X"46",X"43",X"48",X"41",X"61",X"AA",X"B4",X"BA",X"B8",X"BA",X"B7",X"BA",X"AE",X"63",X"49",X"46",
		X"45",X"45",X"46",X"44",X"4D",X"97",X"B6",X"B7",X"BA",X"B7",X"BA",X"B6",X"BB",X"7C",X"4A",X"48",
		X"43",X"46",X"43",X"47",X"42",X"7C",X"B4",X"B5",X"BC",X"B7",X"BC",X"B6",X"BE",X"99",X"52",X"48",
		X"43",X"46",X"43",X"47",X"41",X"60",X"A9",X"B5",X"BA",X"B9",X"BA",X"B8",X"BA",X"B1",X"66",X"47",
		X"45",X"44",X"45",X"45",X"45",X"4A",X"93",X"B7",X"B7",X"BB",X"B8",X"BB",X"B6",X"BC",X"83",X"4B",
		X"47",X"42",X"46",X"43",X"48",X"42",X"75",X"B2",X"B5",X"BC",X"B7",X"BC",X"B6",X"BD",X"A0",X"57",
		X"48",X"43",X"44",X"43",X"46",X"42",X"58",X"A4",X"B6",X"B9",X"BA",X"B9",X"B9",X"B8",X"B6",X"6F",
		X"48",X"46",X"42",X"45",X"43",X"46",X"46",X"88",X"B6",X"B6",X"BC",X"B7",X"BC",X"B5",X"BD",X"90",
		X"4E",X"47",X"42",X"45",X"42",X"47",X"41",X"66",X"AD",X"B5",X"BB",X"B8",X"BA",X"B7",X"BA",X"AD",
		X"62",X"47",X"44",X"43",X"44",X"45",X"45",X"4C",X"95",X"B7",X"B7",X"BB",X"B7",X"BA",X"B4",X"BB",
		X"83",X"4A",X"47",X"42",X"46",X"43",X"48",X"41",X"71",X"B2",X"B5",X"BB",X"B7",X"BA",X"B5",X"BA",
		X"A5",X"5B",X"47",X"44",X"44",X"44",X"46",X"44",X"51",X"9C",X"B7",X"B8",X"BA",X"B7",X"B9",X"B5",
		X"BA",X"7C",X"49",X"47",X"43",X"46",X"43",X"48",X"42",X"77",X"B3",X"B5",X"BC",X"B7",X"BA",X"B5",
		X"BB",X"A2",X"58",X"47",X"44",X"45",X"44",X"47",X"44",X"52",X"9E",X"B7",X"B8",X"BA",X"B7",X"B9",
		X"B4",X"B9",X"7B",X"49",X"47",X"43",X"47",X"44",X"49",X"43",X"76",X"B3",X"B5",X"BB",X"B7",X"BA",
		X"B4",X"BA",X"A4",X"5A",X"47",X"45",X"45",X"45",X"47",X"46",X"51",X"9A",X"B7",X"B7",X"BA",X"B7",
		X"B9",X"B4",X"BA",X"80",X"4A",X"48",X"43",X"47",X"44",X"4A",X"43",X"72",X"B2",X"B5",X"BB",X"B7",
		X"BA",X"B5",X"BA",X"A7",X"5C",X"47",X"45",X"45",X"45",X"47",X"46",X"4F",X"98",X"B7",X"B7",X"BA",
		X"B6",X"BA",X"B4",X"BB",X"84",X"4A",X"48",X"43",X"47",X"44",X"49",X"42",X"6B",X"AF",X"B5",X"BB",
		X"B7",X"B9",X"B6",X"B9",X"AD",X"63",X"48",X"45",X"44",X"45",X"46",X"46",X"4B",X"93",X"B6",X"B6",
		X"BA",X"B6",X"BA",X"B4",X"BC",X"87",X"4C",X"48",X"43",X"47",X"44",X"49",X"41",X"69",X"AE",X"B4",
		X"B9",X"B7",X"B8",X"B6",X"B9",X"AF",X"66",X"48",X"47",X"45",X"46",X"45",X"47",X"47",X"8A",X"B5",
		X"B5",X"BA",X"B5",X"BA",X"B4",X"BD",X"95",X"51",X"49",X"44",X"47",X"44",X"48",X"42",X"5A",X"A5",
		X"B5",X"B8",X"B8",X"B7",X"B8",X"B6",X"B8",X"75",X"49",X"49",X"44",X"47",X"44",X"48",X"42",X"78",
		X"B2",X"B4",X"BA",X"B6",X"BA",X"B5",X"BB",X"A6",X"5B",X"49",X"46",X"46",X"45",X"46",X"44",X"4C",
		X"96",X"B5",X"B6",X"BA",X"B6",X"BA",X"B5",X"BD",X"8A",X"4D",X"49",X"44",X"47",X"43",X"49",X"41",
		X"63",X"AA",X"B4",X"B9",X"B8",X"B9",X"B8",X"B8",X"B5",X"6E",X"48",X"48",X"44",X"47",X"44",X"48",
		X"43",X"7E",X"B3",X"B4",X"BB",X"B6",X"BA",X"B5",X"BC",X"A2",X"59",X"49",X"45",X"46",X"45",X"47",
		X"44",X"4F",X"99",X"B6",X"B7",X"BA",X"B7",X"BA",X"B5",X"BD",X"89",X"4C",X"48",X"43",X"47",X"43",
		X"48",X"41",X"64",X"AB",X"B5",X"BA",X"B8",X"B9",X"B8",X"B8",X"B5",X"6E",X"48",X"47",X"43",X"46",
		X"43",X"47",X"43",X"7E",X"B4",X"B5",X"BB",X"B7",X"BB",X"B6",X"BD",X"A3",X"59",X"48",X"43",X"44",
		X"43",X"45",X"43",X"50",X"9B",X"B6",X"B7",X"BA",X"B8",X"BB",X"B6",X"BC",X"81",X"4A",X"48",X"42",
		X"46",X"42",X"47",X"3F",X"6A",X"AE",X"B5",X"BA",X"B8",X"BA",X"B8",X"B9",X"B2",X"6A",X"48",X"46",
		X"43",X"45",X"43",X"46",X"42",X"80",X"B4",X"B5",X"BB",X"B7",X"BB",X"B6",X"BC",X"A2",X"58",X"48",
		X"44",X"45",X"44",X"45",X"44",X"4C",X"95",X"B6",X"B7",X"BB",X"B7",X"BB",X"B5",X"BD",X"90",X"4E",
		X"48",X"43",X"46",X"43",X"48",X"42",X"5B",X"A5",X"B6",X"B9",X"BA",X"B9",X"BA",X"B6",X"B9",X"7B",
		X"48",X"48",X"42",X"46",X"43",X"49",X"41",X"6E",X"B0",X"B6",X"BB",X"B9",X"BA",X"B8",X"B9",X"B2",
		X"69",X"47",X"46",X"42",X"45",X"43",X"48",X"43",X"7E",X"B5",X"B6",X"BC",X"B8",X"BB",X"B6",X"BC",
		X"A8",X"5D",X"47",X"44",X"44",X"44",X"45",X"46",X"48",X"8E",X"B6",X"B7",X"BC",X"B7",X"BB",X"B5",
		X"BD",X"99",X"52",X"48",X"43",X"45",X"43",X"47",X"44",X"52",X"9D",X"B7",X"B8",X"BB",X"B7",X"BA",
		X"B5",X"BC",X"8A",X"4B",X"48",X"42",X"46",X"43",X"48",X"42",X"5C",X"A6",X"B7",X"B9",X"B9",X"B8",
		X"B9",X"B5",X"B9",X"7C",X"48",X"47",X"41",X"46",X"42",X"49",X"41",X"6A",X"AE",X"B6",X"BA",X"B8",
		X"B9",X"B7",X"B7",X"B3",X"6E",X"46",X"46",X"42",X"46",X"43",X"49",X"41",X"76",X"B3",X"B6",X"BB",
		X"B8",X"BA",X"B6",X"B8",X"AD",X"64",X"46",X"45",X"43",X"46",X"44",X"48",X"45",X"83",X"B5",X"B6",
		X"BB",X"B7",X"BA",X"B5",X"BB",X"A1",X"57",X"47",X"44",X"45",X"45",X"46",X"46",X"4D",X"95",X"B7",
		X"B7",X"BB",X"B7",X"BA",X"B4",X"BC",X"94",X"50",X"48",X"43",X"46",X"44",X"48",X"44",X"54",X"9F",
		X"B7",X"B8",X"BA",X"B7",X"B9",X"B4",X"BB",X"89",X"4C",X"49",X"43",X"47",X"44",X"49",X"43",X"5C",
		X"A6",X"B7",X"B9",X"B9",X"B7",X"B8",X"B4",X"BA",X"82",X"4A",X"49",X"42",X"47",X"43",X"49",X"42",
		X"60",X"A8",X"B6",X"B9",X"B9",X"B7",X"B8",X"B5",X"B9",X"7D",X"49",X"48",X"42",X"47",X"43",X"4A",
		X"41",X"65",X"AB",X"B6",X"B9",X"B8",X"B7",X"B7",X"B5",X"B7",X"78",X"48",X"48",X"43",X"48",X"44",
		X"4A",X"41",X"69",X"AD",X"B5",X"B9",X"B8",X"B8",X"B7",X"B6",X"B6",X"75",X"48",X"48",X"43",X"48",
		X"44",X"4A",X"41",X"6C",X"AF",X"B5",X"B9",X"B7",X"B8",X"B7",X"B7",X"B5",X"71",X"47",X"48",X"43",
		X"48",X"44",X"4A",X"41",X"6F",X"B0",X"B5",X"B9",X"B7",X"B8",X"B7",X"B7",X"B4",X"6F",X"47",X"48",
		X"43",X"48",X"44",X"4A",X"42",X"71",X"B0",X"B5",X"B9",X"B6",X"B8",X"B6",X"B7",X"B3",X"6D",X"47",
		X"48",X"43",X"47",X"44",X"4A",X"42",X"73",X"B1",X"B5",X"BA",X"B7",X"B9",X"B6",X"B8",X"B3",X"6E",
		X"48",X"48",X"43",X"47",X"44",X"49",X"42",X"72",X"B1",X"B4",X"BA",X"B6",X"BA",X"B5",X"BC",X"99",
		X"53",X"49",X"44",X"47",X"43",X"48",X"41",X"67",X"AB",X"B4",X"B9",X"B7",X"B8",X"B7",X"B7",X"B6",
		X"77",X"49",X"49",X"43",X"48",X"43",X"4A",X"40",X"67",X"AC",X"B5",X"B9",X"B8",X"B8",X"B8",X"B7",
		X"B8",X"79",X"49",X"4A",X"43",X"48",X"43",X"4A",X"41",X"65",X"AB",X"B5",X"B9",X"B8",X"B8",X"B9",
		X"B7",X"BA",X"7D",X"4A",X"4A",X"43",X"48",X"43",X"49",X"41",X"61",X"A8",X"B5",X"B8",X"B8",X"B8",
		X"B9",X"B6",X"BB",X"82",X"4B",X"4A",X"43",X"48",X"43",X"49",X"41",X"5D",X"A6",X"B5",X"B8",X"B8",
		X"B7",X"B9",X"B5",X"BB",X"87",X"4C",X"4A",X"43",X"47",X"43",X"48",X"42",X"58",X"A2",X"B5",X"B7",
		X"B9",X"B7",X"B9",X"B5",X"BC",X"8E",X"4E",X"49",X"43",X"47",X"43",X"47",X"42",X"53",X"9D",X"B6",
		X"B7",X"BA",X"B7",X"BA",X"B5",X"BC",X"94",X"50",X"49",X"43",X"46",X"43",X"46",X"43",X"4D",X"95",
		X"B6",X"B6",X"BA",X"B7",X"BA",X"B5",X"BD",X"9C",X"54",X"48",X"43",X"45",X"43",X"46",X"41",X"54",
		X"A0",X"B4",X"B8",X"B9",X"B8",X"B9",X"B7",X"B9",X"7A",X"49",X"49",X"43",X"47",X"43",X"49",X"40",
		X"61",X"A8",X"B5",X"B9",X"B9",X"B8",X"BA",X"B6",X"BB",X"85",X"4B",X"49",X"42",X"46",X"42",X"47",
		X"41",X"56",X"A0",X"B6",X"B7",X"BA",X"B8",X"BB",X"B6",X"BD",X"93",X"4F",X"48",X"43",X"45",X"43",
		X"46",X"44",X"4C",X"95",X"B7",X"B7",X"BB",X"B8",X"BB",X"B6",X"BD",X"A1",X"58",X"48",X"44",X"44",
		X"45",X"44",X"46",X"45",X"87",X"B5",X"B6",X"BB",X"B8",X"BB",X"B7",X"BB",X"AC",X"63",X"47",X"46",
		X"43",X"46",X"43",X"48",X"41",X"78",X"B2",X"B6",X"BB",X"B8",X"BA",X"B8",X"B9",X"B4",X"6D",X"47",
		X"47",X"42",X"46",X"42",X"49",X"40",X"6E",X"AF",X"B6",X"BA",X"B9",X"B9",X"B9",X"B7",X"B8",X"7A",
		X"48",X"48",X"41",X"46",X"42",X"48",X"41",X"5F",X"A7",X"B7",X"B9",X"BA",X"B8",X"BA",X"B5",X"BB",
		X"8A",X"4B",X"48",X"42",X"45",X"43",X"47",X"43",X"51",X"9B",X"B7",X"B8",X"BB",X"B8",X"BA",X"B5",
		X"BC",X"9B",X"53",X"47",X"43",X"44",X"44",X"45",X"46",X"47",X"8A",X"B6",X"B7",X"BB",X"B7",X"BA",
		X"B5",X"BA",X"A9",X"5F",X"46",X"45",X"42",X"46",X"43",X"48",X"41",X"78",X"B3",X"B6",X"BB",X"B8",
		X"B9",X"B7",X"B7",X"B5",X"71",X"45",X"46",X"41",X"46",X"42",X"49",X"40",X"67",X"AC",X"B7",X"BA",
		X"B9",X"B8",X"B9",X"B6",X"B9",X"7F",X"48",X"48",X"42",X"47",X"43",X"48",X"42",X"57",X"A1",X"B7",
		X"B8",X"BB",X"B7",X"B9",X"B4",X"BB",X"97",X"51",X"47",X"43",X"45",X"45",X"46",X"47",X"48",X"8C",
		X"B7",X"B6",X"BB",X"B7",X"BA",X"B5",X"B9",X"AB",X"62",X"46",X"46",X"42",X"47",X"44",X"4A",X"42",
		X"73",X"B1",X"B6",X"BA",X"B8",X"B9",X"B8",X"B6",X"B7",X"7A",X"47",X"48",X"42",X"47",X"43",X"49",
		X"43",X"5A",X"A3",X"B7",X"B8",X"BA",X"B7",X"BA",X"B4",X"BB",X"96",X"51",X"48",X"44",X"46",X"45",
		X"47",X"47",X"49",X"8D",X"B7",X"B6",X"BB",X"B7",X"BA",X"B5",X"B9",X"AB",X"62",X"46",X"47",X"43",
		X"48",X"44",X"4B",X"42",X"71",X"B0",X"B6",X"BA",X"B9",X"B8",X"B8",X"B5",X"B9",X"7F",X"48",X"48",
		X"42",X"47",X"44",X"49",X"44",X"56",X"A0",X"B7",X"B8",X"BA",X"B7",X"B9",X"B4",X"BB",X"9B",X"53",
		X"47",X"44",X"45",X"46",X"46",X"48",X"46",X"87",X"B6",X"B6",X"BB",X"B7",X"B9",X"B6",X"B8",X"B0",
		X"6A",X"46",X"47",X"42",X"48",X"43",X"4A",X"41",X"67",X"AB",X"B6",X"B9",X"B9",X"B7",X"B8",X"B5",
		X"BB",X"89",X"4C",X"49",X"43",X"47",X"44",X"49",X"43",X"56",X"9F",X"B6",X"B7",X"B9",X"B6",X"B9",
		X"B4",X"BB",X"8B",X"4D",X"49",X"43",X"47",X"45",X"48",X"45",X"50",X"98",X"B6",X"B6",X"BA",X"B6",
		X"B9",X"B4",X"BB",X"A4",X"5C",X"48",X"46",X"44",X"47",X"44",X"49",X"42",X"78",X"B2",X"B5",X"B9",
		X"B7",X"B8",X"B7",X"B7",X"B8",X"79",X"48",X"49",X"43",X"48",X"44",X"49",X"42",X"58",X"A1",X"B6",
		X"B6",X"B9",X"B6",X"B9",X"B4",X"BC",X"9B",X"54",X"49",X"45",X"45",X"46",X"45",X"48",X"44",X"82",
		X"B4",X"B5",X"BA",X"B7",X"B9",X"B7",X"B8",X"B4",X"71",X"48",X"49",X"43",X"48",X"43",X"4A",X"41",
		X"60",X"A7",X"B5",X"B7",X"B9",X"B6",X"B9",X"B5",X"BD",X"93",X"50",X"49",X"45",X"46",X"45",X"46",
		X"46",X"47",X"89",X"B5",X"B4",X"B9",X"B6",X"B9",X"B6",X"B9",X"B1",X"6B",X"48",X"49",X"43",X"48",
		X"43",X"4A",X"40",X"63",X"A9",X"B5",X"B8",X"B9",X"B7",X"B9",X"B5",X"BC",X"92",X"50",X"49",X"44",
		X"46",X"45",X"46",X"46",X"47",X"88",X"B5",X"B5",X"BA",X"B7",X"B9",X"B6",X"B9",X"B2",X"6C",X"48",
		X"48",X"42",X"47",X"43",X"49",X"40",X"61",X"A7",X"B5",X"B7",X"B9",X"B7",X"BA",X"B5",X"BD",X"95",
		X"51",X"48",X"44",X"45",X"45",X"45",X"46",X"45",X"85",X"B4",X"B5",X"BA",X"B7",X"BA",X"B7",X"B9",
		X"B3",X"6C",X"46",X"47",X"41",X"46",X"41",X"48",X"3F",X"69",X"AB",X"B6",X"B9",X"B9",X"B8",X"BA",
		X"B7",X"BA",X"82",X"4B",X"48",X"42",X"46",X"42",X"47",X"40",X"6F",X"B0",X"B4",X"BB",X"B7",X"BB",
		X"B6",X"BC",X"A9",X"61",X"48",X"47",X"43",X"46",X"43",X"48",X"40",X"6E",X"AE",X"B5",X"B9",X"B9",
		X"B8",X"B9",X"B7",X"BC",X"8A",X"4D",X"49",X"43",X"46",X"43",X"46",X"44",X"49",X"8F",X"B6",X"B6",
		X"BA",X"B7",X"BA",X"B7",X"BA",X"B0",X"69",X"47",X"48",X"42",X"47",X"42",X"48",X"40",X"61",X"A8",
		X"B6",X"B8",X"BA",X"B7",X"BA",X"B5",X"BD",X"97",X"52",X"49",X"44",X"45",X"45",X"44",X"47",X"43",
		X"80",X"B4",X"B5",X"BA",X"B8",X"B9",X"B8",X"B8",X"B8",X"78",X"48",X"49",X"42",X"47",X"42",X"47",
		X"42",X"53",X"9C",X"B7",X"B7",X"BB",X"B7",X"BB",X"B5",X"BB",X"A7",X"5E",X"46",X"46",X"42",X"46",
		X"42",X"49",X"40",X"6D",X"AE",X"B6",X"B9",X"B9",X"B8",X"B9",X"B5",X"BC",X"8E",X"4D",X"48",X"43",
		X"45",X"44",X"45",X"46",X"47",X"89",X"B6",X"B6",X"BB",X"B8",X"BA",X"B7",X"B8",X"B4",X"72",X"46",
		X"47",X"41",X"46",X"42",X"48",X"41",X"57",X"A0",X"B8",X"B8",X"BB",X"B7",X"BA",X"B5",X"BB",X"A3",
		X"5A",X"46",X"45",X"42",X"46",X"43",X"48",X"40",X"71",X"B0",X"B6",X"BA",X"B9",X"B8",X"B9",X"B5",
		X"BA",X"86",X"4A",X"48",X"42",X"45",X"44",X"46",X"46",X"49",X"8E",X"B7",X"B7",X"BC",X"B8",X"BA",
		X"B6",X"B8",X"B3",X"6F",X"45",X"47",X"41",X"47",X"42",X"49",X"42",X"57",X"A0",X"B8",X"B8",X"BB",
		X"B7",X"BA",X"B5",X"BB",X"A5",X"5C",X"45",X"46",X"43",X"47",X"43",X"4A",X"41",X"6A",X"AD",X"B7",
		X"BA",X"BA",X"B8",X"B9",X"B4",X"BB",X"92",X"4F",X"47",X"44",X"45",X"46",X"45",X"48",X"44",X"80",
		X"B5",X"B6",X"BB",X"B8",X"B9",X"B8",X"B6",X"B8",X"7E",X"48",X"48",X"42",X"47",X"44",X"48",X"46",
		X"4C",X"92",X"B8",X"B7",X"BB",X"B7",X"BA",X"B6",X"B8",X"B1",X"6C",X"46",X"48",X"42",X"48",X"43",
		X"4A",X"43",X"59",X"A2",X"B8",X"B8",X"BB",X"B7",X"BA",X"B4",X"BA",X"A5",X"5C",X"46",X"46",X"43",
		X"48",X"44",X"4B",X"42",X"6A",X"AD",X"B7",X"B9",X"B9",X"B7",X"B9",X"B4",X"BB",X"95",X"50",X"47",
		X"44",X"45",X"46",X"45",X"4A",X"44",X"7C",X"B4",X"B6",X"BA",X"B8",X"B8",X"B8",X"B5",X"BA",X"85",
		X"4A",X"48",X"43",X"47",X"45",X"47",X"47",X"48",X"8A",X"B7",X"B6",X"BB",X"B7",X"B9",X"B6",X"B7",
		X"B6",X"77",X"47",X"48",X"43",X"48",X"44",X"49",X"45",X"50",X"97",X"B7",X"B6",X"BA",X"B5",X"B8",
		X"B4",X"B9",X"AC",X"65",X"46",X"47",X"43",X"48",X"44",X"4B",X"42",X"63",X"A9",X"B7",X"B8",X"B9",
		X"B6",X"B9",X"B4",X"BB",X"9F",X"58",X"47",X"46",X"44",X"47",X"44",X"4A",X"41",X"6D",X"AE",X"B6",
		X"B8",X"B9",X"B6",X"B9",X"B4",X"BC",X"95",X"51",X"48",X"45",X"45",X"47",X"45",X"49",X"43",X"79",
		X"B2",X"B5",X"B9",X"B7",X"B7",X"B7",X"B6",X"B8",X"7B",X"48",X"49",X"43",X"48",X"44",X"49",X"44",
		X"54",X"9C",X"B7",X"B6",X"B9",X"B6",X"B9",X"B5",X"BA",X"AD",X"66",X"47",X"48",X"43",X"48",X"43",
		X"4A",X"42",X"5C",X"A3",X"B7",X"B7",X"BA",X"B6",X"BA",X"B4",X"BB",X"A8",X"60",X"47",X"48",X"44",
		X"48",X"44",X"4A",X"41",X"62",X"A8",X"B6",X"B8",X"B9",X"B7",X"B9",X"B5",X"BA",X"81",X"4A",X"49",
		X"43",X"48",X"43",X"49",X"42",X"5C",X"A4",X"B6",X"B7",X"B9",X"B6",X"B9",X"B4",X"BA",X"A5",X"5D",
		X"47",X"47",X"44",X"48",X"43",X"4A",X"40",X"62",X"A7",X"B6",X"B7",X"B9",X"B6",X"BA",X"B4",X"BB",
		X"A2",X"5B",X"47",X"47",X"44",X"48",X"43",X"4A",X"40",X"65",X"AA",X"B5",X"B8",X"B9",X"B7",X"B9",
		X"B4",X"BC",X"8F",X"4E",X"49",X"44",X"47",X"45",X"47",X"46",X"49",X"8E",X"B6",X"B5",X"BA",X"B7",
		X"B9",X"B7",X"B7",X"B6",X"78",X"47",X"49",X"42",X"47",X"43",X"47",X"44",X"4C",X"90",X"B6",X"B5",
		X"BB",X"B7",X"BA",X"B7",X"B9",X"B6",X"75",X"48",X"49",X"43",X"47",X"44",X"48",X"44",X"4E",X"94",
		X"B7",X"B6",X"BB",X"B7",X"BB",X"B5",X"BD",X"9B",X"54",X"49",X"44",X"46",X"44",X"47",X"45",X"4C",
		X"92",X"B5",X"B5",X"BA",X"B7",X"B9",X"B7",X"B8",X"B5",X"75",X"48",X"49",X"42",X"47",X"43",X"48",
		X"44",X"4C",X"92",X"B6",X"B5",X"BA",X"B6",X"B9",X"B7",X"B8",X"B6",X"76",X"48",X"49",X"43",X"47",
		X"43",X"47",X"44",X"4C",X"92",X"B6",X"B6",X"BB",X"B6",X"BA",X"B5",X"BC",X"A4",X"5A",X"49",X"46",
		X"45",X"46",X"44",X"48",X"43",X"80",X"B3",X"B5",X"BA",X"B8",X"B8",X"B8",X"B6",X"BB",X"89",X"4C",
		X"49",X"43",X"46",X"45",X"45",X"47",X"43",X"7F",X"B4",X"B5",X"BA",X"B8",X"B9",X"B9",X"B6",X"BB",
		X"88",X"4C",X"49",X"44",X"46",X"45",X"45",X"47",X"44",X"7F",X"B4",X"B5",X"BB",X"B7",X"BA",X"B6",
		X"BB",X"A9",X"5F",X"49",X"46",X"45",X"45",X"45",X"47",X"45",X"85",X"B4",X"B5",X"BA",X"B8",X"B9",
		X"B9",X"B7",X"BA",X"86",X"4B",X"49",X"43",X"46",X"44",X"45",X"46",X"43",X"7F",X"B4",X"B5",X"BA",
		X"B9",X"B9",X"BA",X"B6",X"BD",X"8E",X"4E",X"48",X"43",X"44",X"44",X"43",X"47",X"40",X"76",X"B1",
		X"B6",X"B9",X"B9",X"B8",X"BA",X"B6",X"BE",X"97",X"52",X"48",X"45",X"44",X"46",X"43",X"48",X"41",
		X"6D",X"AE",X"B6",X"B9",X"BA",X"B8",X"BB",X"B6",X"BD",X"9F",X"58",X"47",X"46",X"43",X"46",X"42",
		X"49",X"40",X"64",X"A9",X"B7",X"B8",X"BA",X"B7",X"BB",X"B6",X"BC",X"A7",X"5F",X"46",X"47",X"42",
		X"47",X"42",X"49",X"40",X"5A",X"A2",X"B7",X"B7",X"BB",X"B7",X"BB",X"B6",X"BA",X"AD",X"67",X"46",
		X"47",X"41",X"46",X"42",X"48",X"43",X"53",X"9B",X"B8",X"B7",X"BB",X"B8",X"BA",X"B6",X"B8",X"B4",
		X"72",X"46",X"48",X"41",X"46",X"43",X"47",X"44",X"4B",X"90",X"B8",X"B7",X"BB",X"B8",X"BA",X"B8",
		X"B6",X"B8",X"7F",X"48",X"48",X"41",X"45",X"43",X"45",X"46",X"45",X"83",X"B6",X"B7",X"BB",X"B9",
		X"B9",X"B9",X"B5",X"BB",X"8C",X"4C",X"47",X"43",X"44",X"45",X"43",X"48",X"41",X"74",X"B1",X"B7",
		X"BA",X"BA",X"B8",X"BA",X"B4",X"BC",X"9B",X"54",X"46",X"45",X"42",X"46",X"42",X"49",X"40",X"64",
		X"A9",X"B8",X"B9",X"BB",X"B7",X"BA",X"B5",X"BA",X"A9",X"61",X"45",X"47",X"42",X"47",X"42",X"49",
		X"42",X"55",X"9E",X"B8",X"B7",X"BB",X"B7",X"BA",X"B6",X"B8",X"B3",X"70",X"45",X"47",X"41",X"46",
		X"42",X"47",X"43",X"4D",X"94",X"B8",X"B6",X"BB",X"B7",X"B9",X"B6",X"B7",X"B5",X"75",X"46",X"47",
		X"42",X"47",X"44",X"47",X"47",X"48",X"89",X"B7",X"B7",X"BB",X"B8",X"B8",X"B8",X"B5",X"BA",X"8A",
		X"4B",X"47",X"43",X"44",X"46",X"45",X"49",X"42",X"73",X"B1",X"B7",X"B9",X"BA",X"B7",X"B9",X"B4",
		X"BB",X"9F",X"58",X"45",X"46",X"43",X"48",X"44",X"4B",X"42",X"5E",X"A5",X"B8",X"B8",X"BB",X"B7",
		X"BA",X"B4",X"B9",X"AE",X"69",X"45",X"47",X"42",X"48",X"44",X"49",X"45",X"4E",X"93",X"B8",X"B7",
		X"BB",X"B8",X"B9",X"B7",X"B5",X"B8",X"80",X"48",X"48",X"43",X"46",X"46",X"46",X"4A",X"45",X"7C",
		X"B4",X"B7",X"BA",X"B9",X"B8",X"B9",X"B4",X"BB",X"98",X"53",X"47",X"45",X"44",X"47",X"45",X"4B",
		X"43",X"65",X"AA",X"B7",X"B9",X"BA",X"B7",X"BA",X"B4",X"BB",X"8E",X"4D",X"47",X"43",X"45",X"45",
		X"46",X"47",X"4A",X"8E",X"B6",X"B7",X"BA",X"B8",X"B8",X"B7",X"B5",X"B8",X"86",X"49",X"48",X"41",
		X"46",X"44",X"48",X"46",X"4B",X"8E",X"B7",X"B6",X"BC",X"B7",X"BA",X"B6",X"B8",X"B0",X"6B",X"46",
		X"47",X"43",X"47",X"45",X"48",X"47",X"4A",X"8E",X"B7",X"B6",X"BA",X"B8",X"B8",X"B8",X"B6",X"BA",
		X"8A",X"4B",X"49",X"42",X"46",X"43",X"47",X"45",X"4A",X"8D",X"B7",X"B5",X"BB",X"B6",X"B9",X"B5",
		X"B9",X"B1",X"6C",X"46",X"47",X"43",X"47",X"45",X"48",X"47",X"4A",X"8D",X"B7",X"B6",X"BB",X"B8",
		X"B8",X"B8",X"B5",X"BB",X"8B",X"4C",X"48",X"44",X"45",X"47",X"45",X"4A",X"42",X"6F",X"AF",X"B7",
		X"B8",X"B9",X"B6",X"B9",X"B4",X"BB",X"A6",X"5E",X"45",X"47",X"42",X"48",X"43",X"4A",X"43",X"54",
		X"9B",X"B8",X"B6",X"BA",X"B6",X"B9",X"B6",X"B7",X"B7",X"7B",X"48",X"48",X"43",X"47",X"46",X"46",
		X"48",X"44",X"7C",X"B3",X"B6",X"B9",X"B8",X"B7",X"B9",X"B4",X"BC",X"9C",X"56",X"47",X"47",X"44",
		X"48",X"44",X"4B",X"42",X"5C",X"A2",X"B7",X"B6",X"BA",X"B6",X"B9",X"B6",X"B8",X"B4",X"73",X"47",
		X"49",X"43",X"48",X"45",X"47",X"47",X"46",X"83",X"B5",X"B5",X"B9",X"B8",X"B7",X"B9",X"B4",X"BC",
		X"96",X"52",X"47",X"46",X"44",X"48",X"43",X"4A",X"41",X"60",X"A5",X"B6",X"B6",X"BA",X"B6",X"B9",
		X"B5",X"B8",X"B2",X"6F",X"47",X"49",X"43",X"47",X"44",X"47",X"46",X"46",X"86",X"B4",X"B5",X"B9",
		X"B8",X"B8",X"B8",X"B5",X"BC",X"95",X"51",X"48",X"45",X"44",X"47",X"44",X"49",X"41",X"60",X"A6",
		X"B6",X"B7",X"B9",X"B7",X"B9",X"B6",X"B9",X"B0",X"6B",X"46",X"48",X"41",X"47",X"41",X"49",X"3F",
		X"5F",X"A5",X"B6",X"B6",X"BA",X"B6",X"BB",X"B4",X"BD",X"9C",X"57",X"47",X"46",X"44",X"47",X"43",
		X"49",X"41",X"59",X"A1",X"B7",X"B7",X"BA",X"B7",X"B9",X"B7",X"B8",X"B6",X"77",X"47",X"48",X"43",
		X"46",X"44",X"46",X"46",X"44",X"7B",X"B4",X"B4",X"BB",X"B7",X"B9",X"B8",X"B6",X"BA",X"84",X"4A",
		X"48",X"43",X"46",X"44",X"45",X"46",X"46",X"8A",X"B4",X"B7",X"B9",X"B9",X"B8",X"B9",X"B6",X"BB",
		X"92",X"4F",X"49",X"43",X"46",X"43",X"46",X"43",X"51",X"9B",X"B6",X"B7",X"BA",X"B7",X"BB",X"B5",
		X"BE",X"92",X"51",X"48",X"45",X"45",X"46",X"44",X"48",X"41",X"61",X"A9",X"B6",X"B9",X"BA",X"B8",
		X"BA",X"B6",X"BD",X"8E",X"4E",X"49",X"44",X"46",X"45",X"45",X"45",X"49",X"90",X"B5",X"B7",X"B9",
		X"B9",X"B8",X"B9",X"B6",X"BC",X"8F",X"4E",X"4A",X"43",X"46",X"43",X"46",X"43",X"4B",X"91",X"B6",
		X"B5",X"BB",X"B6",X"BB",X"B5",X"BC",X"A6",X"5F",X"47",X"47",X"43",X"46",X"43",X"47",X"43",X"4D",
		X"95",X"B6",X"B7",X"BA",X"B8",X"B8",X"B9",X"B6",X"BC",X"8A",X"4D",X"48",X"44",X"45",X"45",X"44",
		X"48",X"41",X"65",X"AB",X"B6",X"B9",X"B9",X"B8",X"B9",X"B8",X"B9",X"B2",X"6D",X"47",X"49",X"41",
		X"47",X"41",X"48",X"3E",X"60",X"A6",X"B6",X"B7",X"BA",X"B6",X"BB",X"B4",X"BF",X"97",X"55",X"47",
		X"46",X"43",X"47",X"43",X"48",X"40",X"5A",X"A3",X"B7",X"B8",X"BA",X"B8",X"B9",X"B8",X"B8",X"B8",
		X"7A",X"49",X"48",X"44",X"45",X"45",X"44",X"48",X"41",X"75",X"B1",X"B6",X"B9",X"B9",X"B8",X"BA",
		X"B6",X"BB",X"AA",X"62",X"47",X"47",X"43",X"46",X"43",X"46",X"44",X"49",X"8E",X"B6",X"B7",X"BA",
		X"B9",X"B8",X"BA",X"B5",X"BD",X"97",X"52",X"47",X"45",X"43",X"46",X"43",X"48",X"42",X"58",X"A1",
		X"B7",X"B8",X"BA",X"B8",X"B9",X"B8",X"B7",X"BA",X"80",X"4A",X"48",X"44",X"45",X"45",X"44",X"48",
		X"41",X"6E",X"AF",X"B7",X"B9",X"BA",X"B8",X"BA",X"B7",X"BA",X"B0",X"69",X"47",X"47",X"43",X"45",
		X"43",X"46",X"46",X"46",X"86",X"B6",X"B7",X"BA",X"B9",X"B9",X"BA",X"B5",X"BC",X"9F",X"57",X"47",
		X"45",X"43",X"45",X"43",X"47",X"44",X"50",X"99",X"B7",X"B8",X"BA",X"B9",X"B9",X"B9",X"B6",X"BC",
		X"8D",X"4D",X"47",X"43",X"43",X"45",X"43",X"48",X"42",X"5F",X"A7",X"B7",X"B9",X"BB",X"B9",X"B9",
		X"B8",X"B7",X"B7",X"79",X"47",X"47",X"42",X"45",X"44",X"45",X"48",X"43",X"72",X"B2",X"B6",X"BB",
		X"B9",X"B9",X"B9",X"B6",X"BA",X"A7",X"5F",X"44",X"46",X"40",X"46",X"40",X"4A",X"3F",X"5F",X"A4",
		X"B8",X"B7",X"BC",X"B7",X"BB",X"B5",X"BB",X"AB",X"64",X"46",X"46",X"42",X"45",X"44",X"46",X"47",
		X"46",X"88",X"B6",X"B8",X"BA",X"BA",X"B8",X"BA",X"B5",X"BB",X"9F",X"57",X"46",X"44",X"42",X"45",
		X"44",X"47",X"45",X"4F",X"98",X"B7",X"B8",X"BA",X"B9",X"B8",X"B9",X"B5",X"BC",X"91",X"4F",X"46",
		X"43",X"43",X"45",X"44",X"48",X"43",X"58",X"A2",X"B7",X"B9",X"BA",X"B9",X"B8",X"B9",X"B5",X"BA",
		X"83",X"4A",X"47",X"43",X"44",X"45",X"44",X"49",X"42",X"65",X"AC",X"B7",X"BA",X"B9",X"B9",X"B8",
		X"B8",X"B6",X"B7",X"77",X"48",X"47",X"43",X"45",X"45",X"45",X"49",X"43",X"6D",X"B0",X"B6",X"BA",
		X"B8",X"B9",X"B7",X"B7",X"B6",X"B4",X"6F",X"47",X"46",X"43",X"45",X"45",X"46",X"49",X"44",X"76",
		X"B3",X"B5",X"BB",X"B7",X"B9",X"B7",X"B7",X"B6",X"AD",X"64",X"47",X"46",X"43",X"46",X"44",X"49",
		X"43",X"77",X"B2",X"B6",X"BA",X"B8",X"B8",X"B7",X"B6",X"B3",X"6D",X"49",X"46",X"44",X"44",X"46",
		X"45",X"4A",X"43",X"79",X"B2",X"B7",X"BA",X"B9",X"B8",X"B7",X"B6",X"B7",X"AE",X"65",X"48",X"46",
		X"44",X"45",X"46",X"45",X"49",X"45",X"80",X"B5",X"B7",X"BA",X"B8",X"B7",X"B7",X"B4",X"B7",X"A9",
		X"5F",X"47",X"45",X"44",X"45",X"45",X"46",X"48",X"47",X"87",X"B6",X"B7",X"BA",X"B8",X"B7",X"B7",
		X"B4",X"B9",X"A4",X"5A",X"48",X"45",X"45",X"46",X"46",X"47",X"48",X"49",X"8E",X"B6",X"B7",X"BA",
		X"B8",X"B7",X"B7",X"B4",X"BA",X"A0",X"57",X"48",X"45",X"45",X"45",X"46",X"46",X"47",X"4A",X"91",
		X"B6",X"B7",X"B9",X"B8",X"B7",X"B7",X"B4",X"BA",X"9D",X"55",X"48",X"44",X"45",X"46",X"46",X"47",
		X"47",X"4C",X"95",X"B6",X"B8",X"B9",X"B8",X"B6",X"B8",X"B4",X"BB",X"99",X"53",X"48",X"44",X"45",
		X"46",X"46",X"47",X"46",X"4D",X"98",X"B6",X"B8",X"B9",X"B8",X"B7",X"B8",X"B4",X"BB",X"98",X"52",
		X"48",X"44",X"46",X"46",X"47",X"47",X"46",X"4F",X"99",X"B6",X"B8",X"B8",X"B8",X"B6",X"B8",X"B4",
		X"BB",X"97",X"51",X"48",X"45",X"46",X"46",X"47",X"47",X"46",X"4E",X"99",X"B6",X"B8",X"B8",X"B8",
		X"B6",X"B8",X"B4",X"BB",X"96",X"51",X"48",X"44",X"46",X"46",X"46",X"47",X"45",X"4F",X"9A",X"B5",
		X"B7",X"B8",X"B8",X"B6",X"B8",X"B4",X"BB",X"97",X"52",X"49",X"45",X"46",X"46",X"46",X"47",X"45",
		X"4E",X"95",X"B5",X"B6",X"B9",X"B7",X"B8",X"B8",X"B6",X"BA",X"99",X"53",X"49",X"45",X"46",X"47",
		X"44",X"49",X"40",X"6F",X"AD",X"B5",X"B7",X"B9",X"B5",X"BA",X"B3",X"BC",X"97",X"54",X"48",X"46",
		X"45",X"47",X"46",X"47",X"45",X"4D",X"95",X"B5",X"B7",X"B8",X"B8",X"B7",X"B9",X"B5",X"BC",X"9C",
		X"55",X"49",X"45",X"46",X"46",X"46",X"46",X"46",X"49",X"90",X"B5",X"B7",X"BA",X"B9",X"B8",X"B9",
		X"B6",X"BB",X"A3",X"59",X"48",X"45",X"44",X"45",X"45",X"46",X"45",X"48",X"89",X"B6",X"B5",X"BB",
		X"B7",X"BA",X"B8",X"B7",X"B9",X"81",X"4A",X"49",X"43",X"46",X"45",X"45",X"47",X"44",X"84",X"B3",
		X"B7",X"BA",X"B9",X"B9",X"BA",X"B7",X"BB",X"AB",X"61",X"48",X"46",X"44",X"45",X"45",X"45",X"47",
		X"43",X"80",X"B5",X"B6",X"BB",X"B9",X"BA",X"B9",X"B9",X"B9",X"B0",X"64",X"48",X"45",X"44",X"44",
		X"45",X"44",X"48",X"42",X"78",X"B3",X"B6",X"BC",X"B8",X"BB",X"B8",X"BA",X"B7",X"B6",X"6D",X"49",
		X"45",X"44",X"44",X"45",X"44",X"48",X"42",X"6B",X"B0",X"B5",X"BC",X"B8",X"BC",X"B8",X"BB",X"B6",
		X"BA",X"79",X"49",X"46",X"43",X"43",X"44",X"44",X"48",X"42",X"60",X"AA",X"B5",X"BB",X"B9",X"BB",
		X"B7",X"BA",X"B5",X"BC",X"85",X"4B",X"46",X"43",X"44",X"45",X"44",X"47",X"44",X"57",X"A2",X"B7",
		X"B9",X"BA",X"B9",X"B8",X"B8",X"B5",X"B8",X"86",X"4C",X"49",X"44",X"47",X"48",X"48",X"4C",X"46",
		X"6E",X"AA",X"B2",X"B4",X"B4",X"B2",X"B4",X"AF",X"B5",X"9D",X"5F",X"4D",X"4D",X"4B",X"4E",X"4D",
		X"51",X"4E",X"5A",X"97",X"AD",X"AF",X"AF",X"AE",X"AD",X"AD",X"AA",X"AE",X"95",X"5C",X"54",X"50",
		X"52",X"52",X"54",X"54",X"55",X"56",X"8A",X"A8",X"A9",X"AB",X"A9",X"A9",X"A7",X"A7",X"A7",X"9D",
		X"68",X"59",X"56",X"57",X"57",X"59",X"58",X"5C",X"58",X"7D",X"A2",X"A3",X"A6",X"A3",X"A4",X"A2",
		X"A3",X"A0",X"A0",X"74",X"5E",X"5C",X"5C",X"5D",X"5E",X"5E",X"60",X"5E",X"73",X"9A",X"9E",X"A1",
		X"9E",X"9F",X"9D",X"9E",X"9B",X"9E",X"7F",X"64",X"63",X"61",X"62",X"63",X"64",X"65",X"64",X"6D",
		X"91",X"99",X"9B",X"99",X"9A",X"98",X"99",X"96",X"99",X"89",X"6B",X"68",X"66",X"68",X"68",X"69",
		X"69",X"6B",X"6B",X"87",X"94",X"95",X"95",X"94",X"93",X"93",X"92",X"92",X"8D",X"73",X"6D",X"6C",
		X"6D",X"6D",X"6E",X"6E",X"70",X"6F",X"7F",X"8F",X"8F",X"90",X"8E",X"8F",X"8D",X"8D",X"8C",X"8C",
		X"7B",X"72",X"72",X"72",X"73",X"73",X"74",X"75",X"74",X"7A",X"88",X"8A",X"8A",X"89",X"89",X"88",
		X"88",X"87",X"88",X"80",X"78",X"77",X"77",X"78",X"78",X"79",X"7A",X"79",X"7E",X"85",X"85",X"85",
		X"84",X"84",X"83",X"83",X"83",X"81",X"7D",X"7C",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"7F",
		X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"7F",
		X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",
		X"7F",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",
		X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",
		X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",
		X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",
		X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",
		X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",
		X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",
		X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",
		X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",
		X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",
		X"7F",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",
		X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",
		X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",
		X"80",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",X"7F",X"80",
		X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",
		X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",
		X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",
		X"80",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",
		X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",
		X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",
		X"7F",X"7F",X"80",X"80",X"80",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"80",X"80",
		X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"7F",X"80",
		X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F",
		X"80",X"80",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",
		X"80",X"7F",X"7F",X"80",X"80",X"80",X"7F",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"80",X"7F",X"80",X"7F",X"80",X"7F");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
